library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fce0c487",
    12 => x"86c0c84e",
    13 => x"49fce0c4",
    14 => x"48f4c6c4",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087eae9",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"8148731e",
    47 => x"7205a973",
    48 => x"2687f953",
    49 => x"1e731e4f",
    50 => x"c0029a72",
    51 => x"48c087e7",
    52 => x"a9724bc1",
    53 => x"7287d106",
    54 => x"87c90682",
    55 => x"a9728373",
    56 => x"c387f401",
    57 => x"3ab2c187",
    58 => x"8903a972",
    59 => x"c1078073",
    60 => x"f3052b2a",
    61 => x"264b2687",
    62 => x"1e751e4f",
    63 => x"b7714dc4",
    64 => x"b9ff04a1",
    65 => x"bdc381c1",
    66 => x"a2b77207",
    67 => x"c1baff04",
    68 => x"07bdc182",
    69 => x"c187eefe",
    70 => x"b8ff042d",
    71 => x"2d0780c1",
    72 => x"c1b9ff04",
    73 => x"4d260781",
    74 => x"711e4f26",
    75 => x"4966c44a",
    76 => x"c888c148",
    77 => x"997158a6",
    78 => x"1287d402",
    79 => x"08d4ff48",
    80 => x"4966c478",
    81 => x"c888c148",
    82 => x"997158a6",
    83 => x"2687ec05",
    84 => x"4a711e4f",
    85 => x"484966c4",
    86 => x"a6c888c1",
    87 => x"02997158",
    88 => x"d4ff87d6",
    89 => x"78ffc348",
    90 => x"66c45268",
    91 => x"88c14849",
    92 => x"7158a6c8",
    93 => x"87ea0599",
    94 => x"731e4f26",
    95 => x"4bd4ff1e",
    96 => x"6b7bffc3",
    97 => x"7bffc34a",
    98 => x"32c8496b",
    99 => x"ffc3b172",
   100 => x"c84a6b7b",
   101 => x"c3b27131",
   102 => x"496b7bff",
   103 => x"b17232c8",
   104 => x"87c44871",
   105 => x"4c264d26",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4a710e5d",
   109 => x"724cd4ff",
   110 => x"99ffc349",
   111 => x"c6c47c71",
   112 => x"c805bff4",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"ffc329d8",
   117 => x"d07c7199",
   118 => x"29d04966",
   119 => x"7199ffc3",
   120 => x"4966d07c",
   121 => x"ffc329c8",
   122 => x"d07c7199",
   123 => x"ffc34966",
   124 => x"727c7199",
   125 => x"c329d049",
   126 => x"7c7199ff",
   127 => x"f0c94b6c",
   128 => x"ffc34dff",
   129 => x"87d005ab",
   130 => x"6c7cffc3",
   131 => x"028dc14b",
   132 => x"ffc387c6",
   133 => x"87f002ab",
   134 => x"c7fe4873",
   135 => x"49c01e87",
   136 => x"c348d4ff",
   137 => x"81c178ff",
   138 => x"a9b7c8c3",
   139 => x"2687f104",
   140 => x"1e731e4f",
   141 => x"f8c487e7",
   142 => x"1ec04bdf",
   143 => x"c1f0ffc0",
   144 => x"e7fd49f7",
   145 => x"c186c487",
   146 => x"eac005a8",
   147 => x"48d4ff87",
   148 => x"c178ffc3",
   149 => x"c0c0c0c0",
   150 => x"e1c01ec0",
   151 => x"49e9c1f0",
   152 => x"c487c9fd",
   153 => x"05987086",
   154 => x"d4ff87ca",
   155 => x"78ffc348",
   156 => x"87cb48c1",
   157 => x"c187e6fe",
   158 => x"fdfe058b",
   159 => x"fc48c087",
   160 => x"731e87e6",
   161 => x"48d4ff1e",
   162 => x"d378ffc3",
   163 => x"c01ec04b",
   164 => x"c1c1f0ff",
   165 => x"87d4fc49",
   166 => x"987086c4",
   167 => x"ff87ca05",
   168 => x"ffc348d4",
   169 => x"cb48c178",
   170 => x"87f1fd87",
   171 => x"ff058bc1",
   172 => x"48c087db",
   173 => x"0e87f1fb",
   174 => x"0e5c5b5e",
   175 => x"fd4cd4ff",
   176 => x"eac687db",
   177 => x"f0e1c01e",
   178 => x"fb49c8c1",
   179 => x"86c487de",
   180 => x"c802a8c1",
   181 => x"87eafe87",
   182 => x"e2c148c0",
   183 => x"87dafa87",
   184 => x"ffcf4970",
   185 => x"eac699ff",
   186 => x"87c802a9",
   187 => x"c087d3fe",
   188 => x"87cbc148",
   189 => x"c07cffc3",
   190 => x"f4fc4bf1",
   191 => x"02987087",
   192 => x"c087ebc0",
   193 => x"f0ffc01e",
   194 => x"fa49fac1",
   195 => x"86c487de",
   196 => x"d9059870",
   197 => x"7cffc387",
   198 => x"ffc3496c",
   199 => x"7c7c7c7c",
   200 => x"0299c0c1",
   201 => x"48c187c4",
   202 => x"48c087d5",
   203 => x"abc287d1",
   204 => x"c087c405",
   205 => x"c187c848",
   206 => x"fdfe058b",
   207 => x"f948c087",
   208 => x"731e87e4",
   209 => x"f4c6c41e",
   210 => x"c778c148",
   211 => x"48d0ff4b",
   212 => x"c8fb78c2",
   213 => x"48d0ff87",
   214 => x"1ec078c3",
   215 => x"c1d0e5c0",
   216 => x"c7f949c0",
   217 => x"c186c487",
   218 => x"87c105a8",
   219 => x"05abc24b",
   220 => x"48c087c5",
   221 => x"c187f9c0",
   222 => x"d0ff058b",
   223 => x"87f7fc87",
   224 => x"58f8c6c4",
   225 => x"cd059870",
   226 => x"c01ec187",
   227 => x"d0c1f0ff",
   228 => x"87d8f849",
   229 => x"d4ff86c4",
   230 => x"78ffc348",
   231 => x"c487dec4",
   232 => x"ff58fcc6",
   233 => x"78c248d0",
   234 => x"c348d4ff",
   235 => x"48c178ff",
   236 => x"0e87f5f7",
   237 => x"5d5c5b5e",
   238 => x"c34a710e",
   239 => x"d4ff4dff",
   240 => x"ff7c754c",
   241 => x"c3c448d0",
   242 => x"727c7578",
   243 => x"f0ffc01e",
   244 => x"f749d8c1",
   245 => x"86c487d6",
   246 => x"c5029870",
   247 => x"c048c187",
   248 => x"7c7587f0",
   249 => x"c87cfec3",
   250 => x"66d41ec0",
   251 => x"87faf449",
   252 => x"7c7586c4",
   253 => x"7c757c75",
   254 => x"4be0dad8",
   255 => x"496c7c75",
   256 => x"87c50599",
   257 => x"f3058bc1",
   258 => x"ff7c7587",
   259 => x"78c248d0",
   260 => x"cff648c0",
   261 => x"5b5e0e87",
   262 => x"710e5d5c",
   263 => x"c54cc04b",
   264 => x"4adfcdee",
   265 => x"c348d4ff",
   266 => x"496878ff",
   267 => x"05a9fec3",
   268 => x"7087fdc0",
   269 => x"029b734d",
   270 => x"66d087cc",
   271 => x"f449731e",
   272 => x"86c487cf",
   273 => x"d0ff87d6",
   274 => x"78d1c448",
   275 => x"d07dffc3",
   276 => x"88c14866",
   277 => x"7058a6d4",
   278 => x"87f00598",
   279 => x"c348d4ff",
   280 => x"737878ff",
   281 => x"87c5059b",
   282 => x"d048d0ff",
   283 => x"4c4ac178",
   284 => x"fe058ac1",
   285 => x"487487ee",
   286 => x"1e87e9f4",
   287 => x"4a711e73",
   288 => x"d4ff4bc0",
   289 => x"78ffc348",
   290 => x"c448d0ff",
   291 => x"d4ff78c3",
   292 => x"78ffc348",
   293 => x"ffc01e72",
   294 => x"49d1c1f0",
   295 => x"c487cdf4",
   296 => x"05987086",
   297 => x"c0c887d2",
   298 => x"4966cc1e",
   299 => x"c487e6fd",
   300 => x"ff4b7086",
   301 => x"78c248d0",
   302 => x"ebf34873",
   303 => x"5b5e0e87",
   304 => x"c00e5d5c",
   305 => x"f0ffc01e",
   306 => x"f349c9c1",
   307 => x"1ed287de",
   308 => x"49fcc6c4",
   309 => x"c887fefc",
   310 => x"c14cc086",
   311 => x"acb7d284",
   312 => x"c487f804",
   313 => x"bf97fcc6",
   314 => x"99c0c349",
   315 => x"05a9c0c1",
   316 => x"c487e7c0",
   317 => x"bf97c3c7",
   318 => x"c431d049",
   319 => x"bf97c4c7",
   320 => x"7232c84a",
   321 => x"c5c7c4b1",
   322 => x"b14abf97",
   323 => x"ffcf4c71",
   324 => x"c19cffff",
   325 => x"c134ca84",
   326 => x"c7c487e7",
   327 => x"49bf97c5",
   328 => x"99c631c1",
   329 => x"97c6c7c4",
   330 => x"b7c74abf",
   331 => x"c4b1722a",
   332 => x"bf97c1c7",
   333 => x"9dcf4d4a",
   334 => x"97c2c7c4",
   335 => x"9ac34abf",
   336 => x"c7c432ca",
   337 => x"4bbf97c3",
   338 => x"b27333c2",
   339 => x"97c4c7c4",
   340 => x"c0c34bbf",
   341 => x"2bb7c69b",
   342 => x"81c2b273",
   343 => x"307148c1",
   344 => x"48c14970",
   345 => x"4d703075",
   346 => x"84c14c72",
   347 => x"c0c89471",
   348 => x"cc06adb7",
   349 => x"b734c187",
   350 => x"b7c0c82d",
   351 => x"f4ff01ad",
   352 => x"f0487487",
   353 => x"5e0e87de",
   354 => x"0e5d5c5b",
   355 => x"cfc486f8",
   356 => x"78c048e2",
   357 => x"1edac7c4",
   358 => x"defb49c0",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"cec948c0",
   362 => x"c14dc087",
   363 => x"d2fac07e",
   364 => x"c8c449bf",
   365 => x"c8714ad0",
   366 => x"87eeea4b",
   367 => x"c2059870",
   368 => x"c07ec087",
   369 => x"49bfcefa",
   370 => x"4aecc8c4",
   371 => x"ea4bc871",
   372 => x"987087d8",
   373 => x"c087c205",
   374 => x"c0026e7e",
   375 => x"cec487fd",
   376 => x"c44dbfe0",
   377 => x"bf9fd8cf",
   378 => x"d6c5487e",
   379 => x"c705a8ea",
   380 => x"e0cec487",
   381 => x"87ce4dbf",
   382 => x"e9ca486e",
   383 => x"c502a8d5",
   384 => x"c748c087",
   385 => x"c7c487f1",
   386 => x"49751eda",
   387 => x"c487ecf9",
   388 => x"05987086",
   389 => x"48c087c5",
   390 => x"c087dcc7",
   391 => x"49bfcefa",
   392 => x"4aecc8c4",
   393 => x"e94bc871",
   394 => x"987087c0",
   395 => x"c487c805",
   396 => x"c148e2cf",
   397 => x"c087da78",
   398 => x"49bfd2fa",
   399 => x"4ad0c8c4",
   400 => x"e84bc871",
   401 => x"987087e4",
   402 => x"87c5c002",
   403 => x"e6c648c0",
   404 => x"d8cfc487",
   405 => x"c149bf97",
   406 => x"c005a9d5",
   407 => x"cfc487cd",
   408 => x"49bf97d9",
   409 => x"02a9eac2",
   410 => x"c087c5c0",
   411 => x"87c7c648",
   412 => x"97dac7c4",
   413 => x"c3487ebf",
   414 => x"c002a8e9",
   415 => x"486e87ce",
   416 => x"02a8ebc3",
   417 => x"c087c5c0",
   418 => x"87ebc548",
   419 => x"97e5c7c4",
   420 => x"059949bf",
   421 => x"c487ccc0",
   422 => x"bf97e6c7",
   423 => x"02a9c249",
   424 => x"c087c5c0",
   425 => x"87cfc548",
   426 => x"97e7c7c4",
   427 => x"cfc448bf",
   428 => x"4c7058de",
   429 => x"c488c148",
   430 => x"c458e2cf",
   431 => x"bf97e8c7",
   432 => x"c4817549",
   433 => x"bf97e9c7",
   434 => x"7232c84a",
   435 => x"d3c47ea1",
   436 => x"786e48ef",
   437 => x"97eac7c4",
   438 => x"a6c848bf",
   439 => x"e2cfc458",
   440 => x"d4c202bf",
   441 => x"cefac087",
   442 => x"c8c449bf",
   443 => x"c8714aec",
   444 => x"87f6e54b",
   445 => x"c0029870",
   446 => x"48c087c5",
   447 => x"c487f8c3",
   448 => x"4cbfdacf",
   449 => x"5cc3d4c4",
   450 => x"97ffc7c4",
   451 => x"31c849bf",
   452 => x"97fec7c4",
   453 => x"49a14abf",
   454 => x"97c0c8c4",
   455 => x"32d04abf",
   456 => x"c449a172",
   457 => x"bf97c1c8",
   458 => x"7232d84a",
   459 => x"66c449a1",
   460 => x"efd3c491",
   461 => x"d3c481bf",
   462 => x"c8c459f7",
   463 => x"4abf97c7",
   464 => x"c8c432c8",
   465 => x"4bbf97c6",
   466 => x"c8c44aa2",
   467 => x"4bbf97c8",
   468 => x"a27333d0",
   469 => x"c9c8c44a",
   470 => x"cf4bbf97",
   471 => x"7333d89b",
   472 => x"d3c44aa2",
   473 => x"d3c45afb",
   474 => x"c24abff7",
   475 => x"c492748a",
   476 => x"7248fbd3",
   477 => x"cac178a1",
   478 => x"ecc7c487",
   479 => x"c849bf97",
   480 => x"ebc7c431",
   481 => x"a14abf97",
   482 => x"eacfc449",
   483 => x"e6cfc459",
   484 => x"31c549bf",
   485 => x"c981ffc7",
   486 => x"c3d4c429",
   487 => x"f1c7c459",
   488 => x"c84abf97",
   489 => x"f0c7c432",
   490 => x"a24bbf97",
   491 => x"9266c44a",
   492 => x"d3c4826e",
   493 => x"d3c45aff",
   494 => x"78c048f7",
   495 => x"48f3d3c4",
   496 => x"c478a172",
   497 => x"c448c3d4",
   498 => x"78bff7d3",
   499 => x"48c7d4c4",
   500 => x"bffbd3c4",
   501 => x"e2cfc478",
   502 => x"c9c002bf",
   503 => x"c4487487",
   504 => x"c07e7030",
   505 => x"d3c487c9",
   506 => x"c448bfff",
   507 => x"c47e7030",
   508 => x"6e48e6cf",
   509 => x"f848c178",
   510 => x"264d268e",
   511 => x"264b264c",
   512 => x"5b5e0e4f",
   513 => x"710e5d5c",
   514 => x"e2cfc44a",
   515 => x"87cb02bf",
   516 => x"2bc74b72",
   517 => x"ffc14c72",
   518 => x"7287c99c",
   519 => x"722bc84b",
   520 => x"9cffc34c",
   521 => x"bfefd3c4",
   522 => x"cafac083",
   523 => x"d902abbf",
   524 => x"cefac087",
   525 => x"dac7c45b",
   526 => x"f049731e",
   527 => x"86c487fd",
   528 => x"c5059870",
   529 => x"c048c087",
   530 => x"cfc487e6",
   531 => x"d202bfe2",
   532 => x"c4497487",
   533 => x"dac7c491",
   534 => x"cf4d6981",
   535 => x"ffffffff",
   536 => x"7487cb9d",
   537 => x"c491c249",
   538 => x"9f81dac7",
   539 => x"48754d69",
   540 => x"0e87c6fe",
   541 => x"5d5c5b5e",
   542 => x"7186f40e",
   543 => x"c5059c4c",
   544 => x"c348c087",
   545 => x"a4c887f5",
   546 => x"c0486e7e",
   547 => x"0266dc78",
   548 => x"66dc87c7",
   549 => x"c505bf97",
   550 => x"c348c087",
   551 => x"1ec087dd",
   552 => x"c9d049c1",
   553 => x"c886c487",
   554 => x"66c458a6",
   555 => x"87ffc002",
   556 => x"4aeacfc4",
   557 => x"ff4966dc",
   558 => x"7087d4de",
   559 => x"eec00298",
   560 => x"4a66c487",
   561 => x"cb4966dc",
   562 => x"f7deff4b",
   563 => x"02987087",
   564 => x"1ec087dd",
   565 => x"c40266c8",
   566 => x"c24dc087",
   567 => x"754dc187",
   568 => x"87cacf49",
   569 => x"a6c886c4",
   570 => x"0566c458",
   571 => x"c487c1ff",
   572 => x"c4c20266",
   573 => x"81dc4987",
   574 => x"7869486e",
   575 => x"da4966c4",
   576 => x"4da4c481",
   577 => x"c47d699f",
   578 => x"02bfe2cf",
   579 => x"66c487d5",
   580 => x"9f81d449",
   581 => x"ffc04969",
   582 => x"487199ff",
   583 => x"a6cc30d0",
   584 => x"c887c558",
   585 => x"78c048a6",
   586 => x"484966c8",
   587 => x"7d70806d",
   588 => x"a4cc7cc0",
   589 => x"d0796d49",
   590 => x"79c049a4",
   591 => x"c048a6c4",
   592 => x"4aa4d478",
   593 => x"c84966c4",
   594 => x"49a17291",
   595 => x"796d41c0",
   596 => x"c14866c4",
   597 => x"58a6c880",
   598 => x"04a8b7c6",
   599 => x"6e87e2ff",
   600 => x"2ac94abf",
   601 => x"f0c04972",
   602 => x"d8ddff4a",
   603 => x"c14a7087",
   604 => x"7249a4c4",
   605 => x"c248c179",
   606 => x"f448c087",
   607 => x"87f9f98e",
   608 => x"5c5b5e0e",
   609 => x"4c710e5d",
   610 => x"cac1029c",
   611 => x"49a4c887",
   612 => x"c2c10269",
   613 => x"4a66d087",
   614 => x"d482496c",
   615 => x"66d05aa6",
   616 => x"cfc4b94d",
   617 => x"ff4abfde",
   618 => x"719972ba",
   619 => x"e4c00299",
   620 => x"4ba4c487",
   621 => x"c8f9496b",
   622 => x"c47b7087",
   623 => x"49bfdacf",
   624 => x"7c71816c",
   625 => x"cfc4b975",
   626 => x"ff4abfde",
   627 => x"719972ba",
   628 => x"dcff0599",
   629 => x"f87c7587",
   630 => x"731e87df",
   631 => x"9b4b711e",
   632 => x"c887c702",
   633 => x"056949a3",
   634 => x"48c087c5",
   635 => x"c487f7c0",
   636 => x"4abff3d3",
   637 => x"6949a3c4",
   638 => x"c489c249",
   639 => x"91bfdacf",
   640 => x"c44aa271",
   641 => x"49bfdecf",
   642 => x"a271996b",
   643 => x"cefac04a",
   644 => x"1e66c85a",
   645 => x"e2e94972",
   646 => x"7086c487",
   647 => x"87c40598",
   648 => x"87c248c0",
   649 => x"d4f748c1",
   650 => x"1e731e87",
   651 => x"029b4b71",
   652 => x"a3c887c7",
   653 => x"c5056949",
   654 => x"c048c087",
   655 => x"d3c487f7",
   656 => x"c44abff3",
   657 => x"496949a3",
   658 => x"cfc489c2",
   659 => x"7191bfda",
   660 => x"cfc44aa2",
   661 => x"6b49bfde",
   662 => x"4aa27199",
   663 => x"5acefac0",
   664 => x"721e66c8",
   665 => x"87cbe549",
   666 => x"987086c4",
   667 => x"c087c405",
   668 => x"c187c248",
   669 => x"87c5f648",
   670 => x"5c5b5e0e",
   671 => x"86f80e5d",
   672 => x"7eff4c71",
   673 => x"6949a4c8",
   674 => x"d44bc04d",
   675 => x"49734aa4",
   676 => x"a17291c8",
   677 => x"d8496949",
   678 => x"8a714a66",
   679 => x"d85aa6c8",
   680 => x"cc01a966",
   681 => x"b766c487",
   682 => x"87c506ad",
   683 => x"66c47e73",
   684 => x"c683c14d",
   685 => x"ff04abb7",
   686 => x"486e87d1",
   687 => x"f8f48ef8",
   688 => x"5b5e0e87",
   689 => x"f00e5d5c",
   690 => x"6e7e7186",
   691 => x"c481c849",
   692 => x"786948a6",
   693 => x"78ff80c4",
   694 => x"a6d04dc0",
   695 => x"6e4cc05d",
   696 => x"7483d44b",
   697 => x"7392c84a",
   698 => x"66cc4aa2",
   699 => x"7391c849",
   700 => x"486a49a1",
   701 => x"49708869",
   702 => x"adb7c04d",
   703 => x"0d87c203",
   704 => x"ac66cc8d",
   705 => x"c487cd02",
   706 => x"03adb766",
   707 => x"a6cc87c6",
   708 => x"5da6c85c",
   709 => x"b7c684c1",
   710 => x"c2ff04ac",
   711 => x"4866cc87",
   712 => x"a6d080c1",
   713 => x"a8b7c658",
   714 => x"87f1fe04",
   715 => x"f04866c8",
   716 => x"87c5f38e",
   717 => x"5c5b5e0e",
   718 => x"86f00e5d",
   719 => x"e0c04b71",
   720 => x"28c94866",
   721 => x"7358a6c8",
   722 => x"c6c3029b",
   723 => x"49a3c887",
   724 => x"fec20269",
   725 => x"decfc487",
   726 => x"b9ff49bf",
   727 => x"66c44871",
   728 => x"58a6cc98",
   729 => x"9d6b4d71",
   730 => x"6c4ca3c4",
   731 => x"ad66c87e",
   732 => x"c487c605",
   733 => x"c8c27b66",
   734 => x"1e66c887",
   735 => x"f7fb4973",
   736 => x"d086c487",
   737 => x"b7c058a6",
   738 => x"87d104a8",
   739 => x"cc4aa3d4",
   740 => x"91c84966",
   741 => x"2149a172",
   742 => x"c77c697b",
   743 => x"cc7bc087",
   744 => x"7c6949a3",
   745 => x"6b4866c4",
   746 => x"58a6c888",
   747 => x"49731e75",
   748 => x"c487c5fb",
   749 => x"58a6d086",
   750 => x"49a3c4c1",
   751 => x"06ad4a69",
   752 => x"cc87f3c0",
   753 => x"b7c04866",
   754 => x"e9c004a8",
   755 => x"48a6c887",
   756 => x"cc78a3d4",
   757 => x"91c84966",
   758 => x"758166c8",
   759 => x"70886948",
   760 => x"06a97249",
   761 => x"497387d0",
   762 => x"7087d6fb",
   763 => x"c891c849",
   764 => x"41758166",
   765 => x"66c4796e",
   766 => x"49731e49",
   767 => x"c487c1f6",
   768 => x"dac7c486",
   769 => x"f749731e",
   770 => x"86c487d0",
   771 => x"c049a3d0",
   772 => x"f07966e0",
   773 => x"87e1ef8e",
   774 => x"711e731e",
   775 => x"c0029b4b",
   776 => x"d4c487e4",
   777 => x"4a735bc7",
   778 => x"cfc48ac2",
   779 => x"9249bfda",
   780 => x"bff3d3c4",
   781 => x"c4807248",
   782 => x"7158cbd4",
   783 => x"c430c448",
   784 => x"c058eacf",
   785 => x"d4c487ed",
   786 => x"d3c448c3",
   787 => x"c478bff7",
   788 => x"c448c7d4",
   789 => x"78bffbd3",
   790 => x"bfe2cfc4",
   791 => x"c487c902",
   792 => x"49bfdacf",
   793 => x"87c731c4",
   794 => x"bfffd3c4",
   795 => x"c431c449",
   796 => x"ee59eacf",
   797 => x"5e0e87c7",
   798 => x"710e5c5b",
   799 => x"724bc04a",
   800 => x"e1c0029a",
   801 => x"49a2da87",
   802 => x"c44b699f",
   803 => x"02bfe2cf",
   804 => x"a2d487cf",
   805 => x"49699f49",
   806 => x"ffffc04c",
   807 => x"c234d09c",
   808 => x"744cc087",
   809 => x"4973b349",
   810 => x"ed87edfd",
   811 => x"5e0e87cd",
   812 => x"0e5d5c5b",
   813 => x"4a7186f4",
   814 => x"9a727ec0",
   815 => x"c487d802",
   816 => x"c048d6c7",
   817 => x"cec7c478",
   818 => x"c7d4c448",
   819 => x"c7c478bf",
   820 => x"d4c448d2",
   821 => x"c478bfc3",
   822 => x"c048f7cf",
   823 => x"e6cfc450",
   824 => x"c7c449bf",
   825 => x"714abfd6",
   826 => x"cac403aa",
   827 => x"cf497287",
   828 => x"eac00599",
   829 => x"cafac087",
   830 => x"cec7c448",
   831 => x"c7c478bf",
   832 => x"c7c41eda",
   833 => x"c449bfce",
   834 => x"c148cec7",
   835 => x"ff7178a1",
   836 => x"c487e8dd",
   837 => x"c6fac086",
   838 => x"dac7c448",
   839 => x"c087cc78",
   840 => x"48bfc6fa",
   841 => x"c080e0c0",
   842 => x"c458cafa",
   843 => x"48bfd6c7",
   844 => x"c7c480c1",
   845 => x"862758da",
   846 => x"bf00000e",
   847 => x"9d4dbf97",
   848 => x"87e3c202",
   849 => x"02ade5c3",
   850 => x"c087dcc2",
   851 => x"4bbfc6fa",
   852 => x"1149a3cb",
   853 => x"05accf4c",
   854 => x"7587d2c1",
   855 => x"c199df49",
   856 => x"c491cd89",
   857 => x"c181eacf",
   858 => x"51124aa3",
   859 => x"124aa3c3",
   860 => x"4aa3c551",
   861 => x"a3c75112",
   862 => x"c951124a",
   863 => x"51124aa3",
   864 => x"124aa3ce",
   865 => x"4aa3d051",
   866 => x"a3d25112",
   867 => x"d451124a",
   868 => x"51124aa3",
   869 => x"124aa3d6",
   870 => x"4aa3d851",
   871 => x"a3dc5112",
   872 => x"de51124a",
   873 => x"51124aa3",
   874 => x"fac07ec1",
   875 => x"c8497487",
   876 => x"ebc00599",
   877 => x"d0497487",
   878 => x"87d10599",
   879 => x"c00266dc",
   880 => x"497387cb",
   881 => x"700f66dc",
   882 => x"d3c00298",
   883 => x"c0056e87",
   884 => x"cfc487c6",
   885 => x"50c048ea",
   886 => x"bfc6fac0",
   887 => x"87e1c248",
   888 => x"48f7cfc4",
   889 => x"c47e50c0",
   890 => x"49bfe6cf",
   891 => x"bfd6c7c4",
   892 => x"04aa714a",
   893 => x"c487f6fb",
   894 => x"05bfc7d4",
   895 => x"c487c8c0",
   896 => x"02bfe2cf",
   897 => x"c487f8c1",
   898 => x"49bfd2c7",
   899 => x"7087f2e7",
   900 => x"d6c7c449",
   901 => x"48a6c459",
   902 => x"bfd2c7c4",
   903 => x"e2cfc478",
   904 => x"d8c002bf",
   905 => x"4966c487",
   906 => x"ffffffcf",
   907 => x"02a999f8",
   908 => x"c087c5c0",
   909 => x"87e1c04c",
   910 => x"dcc04cc1",
   911 => x"4966c487",
   912 => x"99f8ffcf",
   913 => x"c8c002a9",
   914 => x"48a6c887",
   915 => x"c5c078c0",
   916 => x"48a6c887",
   917 => x"66c878c1",
   918 => x"059c744c",
   919 => x"c487e0c0",
   920 => x"89c24966",
   921 => x"bfdacfc4",
   922 => x"d3c4914a",
   923 => x"c44abff3",
   924 => x"7248cec7",
   925 => x"c7c478a1",
   926 => x"78c048d6",
   927 => x"c087def9",
   928 => x"e58ef448",
   929 => x"000087f3",
   930 => x"ffff0000",
   931 => x"0e96ffff",
   932 => x"0e9f0000",
   933 => x"41460000",
   934 => x"20323354",
   935 => x"46002020",
   936 => x"36315441",
   937 => x"00202020",
   938 => x"48d0ff1e",
   939 => x"2678e0c0",
   940 => x"f8c21e4f",
   941 => x"497087cd",
   942 => x"87c60299",
   943 => x"05a9fbc0",
   944 => x"487187f0",
   945 => x"5e0e4f26",
   946 => x"710e5c5b",
   947 => x"c24cc04b",
   948 => x"7087f0f7",
   949 => x"c0029949",
   950 => x"ecc087fa",
   951 => x"f3c002a9",
   952 => x"a9fbc087",
   953 => x"87ecc002",
   954 => x"acb766cc",
   955 => x"d087c703",
   956 => x"87c20266",
   957 => x"99715371",
   958 => x"c187c202",
   959 => x"c2f7c284",
   960 => x"99497087",
   961 => x"c087cd02",
   962 => x"c702a9ec",
   963 => x"a9fbc087",
   964 => x"87d4ff05",
   965 => x"c30266d0",
   966 => x"7b97c087",
   967 => x"05a9ecc0",
   968 => x"4a7487c4",
   969 => x"4a7487c5",
   970 => x"728a0ac0",
   971 => x"2687c248",
   972 => x"264c264d",
   973 => x"1e4f264b",
   974 => x"87c7f6c2",
   975 => x"c04a4970",
   976 => x"c904aaf0",
   977 => x"aaf9c087",
   978 => x"c087c301",
   979 => x"c1c18af0",
   980 => x"87c904aa",
   981 => x"01aadac1",
   982 => x"f7c087c3",
   983 => x"2648728a",
   984 => x"5b5e0e4f",
   985 => x"4a710e5c",
   986 => x"724cd4ff",
   987 => x"87e9c049",
   988 => x"029b4b70",
   989 => x"8bc187c2",
   990 => x"c548d0ff",
   991 => x"7cd5c178",
   992 => x"31c64973",
   993 => x"97cdebc1",
   994 => x"71484abf",
   995 => x"ff7c70b0",
   996 => x"78c448d0",
   997 => x"d8fe4873",
   998 => x"5b5e0e87",
   999 => x"f80e5d5c",
  1000 => x"c04c7186",
  1001 => x"fdf4c27e",
  1002 => x"c14bc087",
  1003 => x"bf97cbc1",
  1004 => x"04a9c049",
  1005 => x"f8fb87cf",
  1006 => x"c183c187",
  1007 => x"bf97cbc1",
  1008 => x"f106ab49",
  1009 => x"cbc1c187",
  1010 => x"d002bf97",
  1011 => x"f2f3c287",
  1012 => x"99497087",
  1013 => x"c087c602",
  1014 => x"f005a9ec",
  1015 => x"c24bc087",
  1016 => x"7087e0f3",
  1017 => x"daf3c24d",
  1018 => x"58a6c887",
  1019 => x"87d3f3c2",
  1020 => x"83c14a70",
  1021 => x"9749a4c8",
  1022 => x"02ad4969",
  1023 => x"ffc087c7",
  1024 => x"e7c005ad",
  1025 => x"49a4c987",
  1026 => x"c4496997",
  1027 => x"c702a966",
  1028 => x"ffc04887",
  1029 => x"87d405a8",
  1030 => x"9749a4ca",
  1031 => x"02aa4969",
  1032 => x"ffc087c6",
  1033 => x"87c405aa",
  1034 => x"87d07ec1",
  1035 => x"02adecc0",
  1036 => x"fbc087c6",
  1037 => x"87c405ad",
  1038 => x"7ec14bc0",
  1039 => x"defe026e",
  1040 => x"87e4f987",
  1041 => x"8ef84873",
  1042 => x"0087e4fb",
  1043 => x"5c5b5e0e",
  1044 => x"86f80e5d",
  1045 => x"d4ff4d71",
  1046 => x"c41e754b",
  1047 => x"e049d0d4",
  1048 => x"86c487d1",
  1049 => x"c4029870",
  1050 => x"a6c487cc",
  1051 => x"cfebc148",
  1052 => x"497578bf",
  1053 => x"ff87eafb",
  1054 => x"78c548d0",
  1055 => x"c07bd6c1",
  1056 => x"49a2754a",
  1057 => x"82c17b11",
  1058 => x"04aab7cb",
  1059 => x"4acc87f3",
  1060 => x"c17bffc3",
  1061 => x"b7e0c082",
  1062 => x"87f404aa",
  1063 => x"c448d0ff",
  1064 => x"7bffc378",
  1065 => x"d3c178c5",
  1066 => x"c47bc17b",
  1067 => x"c0486678",
  1068 => x"c206a8b7",
  1069 => x"d4c487f0",
  1070 => x"c44cbfd8",
  1071 => x"88744866",
  1072 => x"7458a6c8",
  1073 => x"f9c1029c",
  1074 => x"dac7c487",
  1075 => x"4dc0c87e",
  1076 => x"acb7c08c",
  1077 => x"c887c603",
  1078 => x"c04da4c0",
  1079 => x"cbd4c44c",
  1080 => x"d049bf97",
  1081 => x"87d10299",
  1082 => x"d4c41ec0",
  1083 => x"e9e349d0",
  1084 => x"7086c487",
  1085 => x"eec04a49",
  1086 => x"dac7c487",
  1087 => x"d0d4c41e",
  1088 => x"87d6e349",
  1089 => x"497086c4",
  1090 => x"48d0ff4a",
  1091 => x"c178c5c8",
  1092 => x"976e7bd4",
  1093 => x"486e7bbf",
  1094 => x"7e7080c1",
  1095 => x"ff058dc1",
  1096 => x"d0ff87f0",
  1097 => x"7278c448",
  1098 => x"87c5059a",
  1099 => x"c7c148c0",
  1100 => x"c41ec187",
  1101 => x"e149d0d4",
  1102 => x"86c487c6",
  1103 => x"fe059c74",
  1104 => x"66c487c7",
  1105 => x"a8b7c048",
  1106 => x"c487d106",
  1107 => x"c048d0d4",
  1108 => x"c080d078",
  1109 => x"c480f478",
  1110 => x"78bfdcd4",
  1111 => x"c04866c4",
  1112 => x"fd01a8b7",
  1113 => x"d0ff87d0",
  1114 => x"c178c548",
  1115 => x"7bc07bd3",
  1116 => x"48c178c4",
  1117 => x"48c087c2",
  1118 => x"4d268ef8",
  1119 => x"4b264c26",
  1120 => x"5e0e4f26",
  1121 => x"0e5d5c5b",
  1122 => x"c04b711e",
  1123 => x"04ab4d4c",
  1124 => x"c087e8c0",
  1125 => x"751ed9fe",
  1126 => x"87c4029d",
  1127 => x"87c24ac0",
  1128 => x"49724ac1",
  1129 => x"c487c7ec",
  1130 => x"c17e7086",
  1131 => x"c2056e84",
  1132 => x"c14c7387",
  1133 => x"06ac7385",
  1134 => x"6e87d8ff",
  1135 => x"f9fe2648",
  1136 => x"5b5e0e87",
  1137 => x"1e0e5d5c",
  1138 => x"de494c71",
  1139 => x"ecd5c491",
  1140 => x"9785714d",
  1141 => x"ddc1026d",
  1142 => x"d8d5c487",
  1143 => x"82744abf",
  1144 => x"ddfe4972",
  1145 => x"6e7e7087",
  1146 => x"87f3c002",
  1147 => x"4be0d5c4",
  1148 => x"49cb4a6e",
  1149 => x"87f0fafe",
  1150 => x"93cb4b74",
  1151 => x"83e1ebc1",
  1152 => x"c8c183c4",
  1153 => x"49747bfa",
  1154 => x"87cbcfc1",
  1155 => x"ebc17b75",
  1156 => x"49bf97ce",
  1157 => x"e0d5c41e",
  1158 => x"d9eec249",
  1159 => x"7486c487",
  1160 => x"f2cec149",
  1161 => x"c149c087",
  1162 => x"c487d1d0",
  1163 => x"c048ccd4",
  1164 => x"dd49c178",
  1165 => x"fd2687e1",
  1166 => x"6f4c87c0",
  1167 => x"6e696461",
  1168 => x"2e2e2e67",
  1169 => x"5b5e0e00",
  1170 => x"4b710e5c",
  1171 => x"d8d5c44a",
  1172 => x"497282bf",
  1173 => x"7087ebfc",
  1174 => x"c4029c4c",
  1175 => x"d5e84987",
  1176 => x"d8d5c487",
  1177 => x"c178c048",
  1178 => x"87ebdc49",
  1179 => x"0e87cdfc",
  1180 => x"5d5c5b5e",
  1181 => x"c486f40e",
  1182 => x"c04ddac7",
  1183 => x"48a6c44c",
  1184 => x"d5c478c0",
  1185 => x"c049bfd8",
  1186 => x"c1c106a9",
  1187 => x"dac7c487",
  1188 => x"c0029848",
  1189 => x"fec087f8",
  1190 => x"66c81ed9",
  1191 => x"c487c702",
  1192 => x"78c048a6",
  1193 => x"a6c487c5",
  1194 => x"c478c148",
  1195 => x"fde74966",
  1196 => x"7086c487",
  1197 => x"c484c14d",
  1198 => x"80c14866",
  1199 => x"c458a6c8",
  1200 => x"49bfd8d5",
  1201 => x"87c603ac",
  1202 => x"ff059d75",
  1203 => x"4cc087c8",
  1204 => x"c3029d75",
  1205 => x"fec087e0",
  1206 => x"66c81ed9",
  1207 => x"cc87c702",
  1208 => x"78c048a6",
  1209 => x"a6cc87c5",
  1210 => x"cc78c148",
  1211 => x"fde64966",
  1212 => x"7086c487",
  1213 => x"c2026e7e",
  1214 => x"496e87e9",
  1215 => x"699781cb",
  1216 => x"0299d049",
  1217 => x"c187d6c1",
  1218 => x"744ac5c9",
  1219 => x"c191cb49",
  1220 => x"7281e1eb",
  1221 => x"c381c879",
  1222 => x"497451ff",
  1223 => x"d5c491de",
  1224 => x"85714dec",
  1225 => x"7d97c1c2",
  1226 => x"c049a5c1",
  1227 => x"cfc451e0",
  1228 => x"02bf97ea",
  1229 => x"84c187d2",
  1230 => x"c44ba5c2",
  1231 => x"db4aeacf",
  1232 => x"e3f5fe49",
  1233 => x"87dbc187",
  1234 => x"c049a5cd",
  1235 => x"c284c151",
  1236 => x"4a6e4ba5",
  1237 => x"f5fe49cb",
  1238 => x"c6c187ce",
  1239 => x"c1c7c187",
  1240 => x"cb49744a",
  1241 => x"e1ebc191",
  1242 => x"c4797281",
  1243 => x"bf97eacf",
  1244 => x"7487d802",
  1245 => x"c191de49",
  1246 => x"ecd5c484",
  1247 => x"c483714b",
  1248 => x"dd4aeacf",
  1249 => x"dff4fe49",
  1250 => x"7487d887",
  1251 => x"c493de4b",
  1252 => x"cb83ecd5",
  1253 => x"51c049a3",
  1254 => x"6e7384c1",
  1255 => x"fe49cb4a",
  1256 => x"c487c5f4",
  1257 => x"80c14866",
  1258 => x"c758a6c8",
  1259 => x"c5c003ac",
  1260 => x"fc056e87",
  1261 => x"487487e0",
  1262 => x"fdf68ef4",
  1263 => x"1e731e87",
  1264 => x"cb494b71",
  1265 => x"e1ebc191",
  1266 => x"4aa1c881",
  1267 => x"48cdebc1",
  1268 => x"a1c95012",
  1269 => x"cbc1c14a",
  1270 => x"ca501248",
  1271 => x"ceebc181",
  1272 => x"c1501148",
  1273 => x"bf97ceeb",
  1274 => x"49c01e49",
  1275 => x"87c6e7c2",
  1276 => x"48ccd4c4",
  1277 => x"49c178de",
  1278 => x"2687dcd6",
  1279 => x"1e87fff5",
  1280 => x"cb494a71",
  1281 => x"e1ebc191",
  1282 => x"1181c881",
  1283 => x"d0d4c448",
  1284 => x"d8d5c458",
  1285 => x"c178c048",
  1286 => x"87fbd549",
  1287 => x"c01e4f26",
  1288 => x"d7c8c149",
  1289 => x"1e4f2687",
  1290 => x"d2029971",
  1291 => x"f6ecc187",
  1292 => x"f750c048",
  1293 => x"ffcfc180",
  1294 => x"daebc140",
  1295 => x"c187ce78",
  1296 => x"c148f2ec",
  1297 => x"fc78d3eb",
  1298 => x"ded0c180",
  1299 => x"0e4f2678",
  1300 => x"0e5c5b5e",
  1301 => x"cb4a4c71",
  1302 => x"e1ebc192",
  1303 => x"49a2c882",
  1304 => x"974ba2c9",
  1305 => x"971e4b6b",
  1306 => x"ca1e4969",
  1307 => x"c0491282",
  1308 => x"c087d1f3",
  1309 => x"87dfd449",
  1310 => x"c5c14974",
  1311 => x"8ef887d9",
  1312 => x"1e87f9f3",
  1313 => x"4b711e73",
  1314 => x"87c3ff49",
  1315 => x"fefe4973",
  1316 => x"87eaf387",
  1317 => x"711e731e",
  1318 => x"4aa3c64b",
  1319 => x"c187db02",
  1320 => x"87d6028a",
  1321 => x"dac1028a",
  1322 => x"c0028a87",
  1323 => x"028a87fc",
  1324 => x"8a87e1c0",
  1325 => x"c187cb02",
  1326 => x"49c787db",
  1327 => x"c187c0fd",
  1328 => x"d5c487de",
  1329 => x"c102bfd8",
  1330 => x"c14887cb",
  1331 => x"dcd5c488",
  1332 => x"87c1c158",
  1333 => x"bfdcd5c4",
  1334 => x"87f9c002",
  1335 => x"bfd8d5c4",
  1336 => x"c480c148",
  1337 => x"c058dcd5",
  1338 => x"d5c487eb",
  1339 => x"c649bfd8",
  1340 => x"dcd5c489",
  1341 => x"a9b7c059",
  1342 => x"c487da03",
  1343 => x"c048d8d5",
  1344 => x"c487d278",
  1345 => x"02bfdcd5",
  1346 => x"d5c487cb",
  1347 => x"c648bfd8",
  1348 => x"dcd5c480",
  1349 => x"d149c058",
  1350 => x"497387fd",
  1351 => x"87f7c2c1",
  1352 => x"0e87dbf1",
  1353 => x"5d5c5b5e",
  1354 => x"86d0ff0e",
  1355 => x"c859a6dc",
  1356 => x"78c048a6",
  1357 => x"c4c180c4",
  1358 => x"80c47866",
  1359 => x"80c478c1",
  1360 => x"d5c478c1",
  1361 => x"78c148dc",
  1362 => x"bfccd4c4",
  1363 => x"05a8de48",
  1364 => x"daf487cb",
  1365 => x"cc497087",
  1366 => x"f9cf59a6",
  1367 => x"c5dec287",
  1368 => x"87cde587",
  1369 => x"87dbddc2",
  1370 => x"fbc04c70",
  1371 => x"fbc102ac",
  1372 => x"0566d887",
  1373 => x"c187edc1",
  1374 => x"c44a66c0",
  1375 => x"727e6a82",
  1376 => x"cbe6c11e",
  1377 => x"4966c448",
  1378 => x"204aa1c8",
  1379 => x"05aa7141",
  1380 => x"511087f9",
  1381 => x"c0c14a26",
  1382 => x"cec14866",
  1383 => x"496a78fd",
  1384 => x"517481c7",
  1385 => x"4966c0c1",
  1386 => x"51c181c8",
  1387 => x"4966c0c1",
  1388 => x"51c081c9",
  1389 => x"4966c0c1",
  1390 => x"51c081ca",
  1391 => x"1ed81ec1",
  1392 => x"81c8496a",
  1393 => x"c887ffe3",
  1394 => x"66c4c186",
  1395 => x"01a8c048",
  1396 => x"a6c887c7",
  1397 => x"ce78c148",
  1398 => x"66c4c187",
  1399 => x"d088c148",
  1400 => x"87c358a6",
  1401 => x"d087cae3",
  1402 => x"78c248a6",
  1403 => x"cd029c74",
  1404 => x"66c887e0",
  1405 => x"66c8c148",
  1406 => x"d5cd03a8",
  1407 => x"48a6dc87",
  1408 => x"80e878c0",
  1409 => x"dac278c0",
  1410 => x"4c7087f9",
  1411 => x"05acd0c1",
  1412 => x"c487dac2",
  1413 => x"dee47e66",
  1414 => x"c8497087",
  1415 => x"dac259a6",
  1416 => x"4c7087e1",
  1417 => x"05acecc0",
  1418 => x"c887edc1",
  1419 => x"91cb4966",
  1420 => x"8166c0c1",
  1421 => x"6a4aa1c4",
  1422 => x"4aa1c84d",
  1423 => x"c15266c4",
  1424 => x"c279ffcf",
  1425 => x"7087fcd9",
  1426 => x"d9029c4c",
  1427 => x"acfbc087",
  1428 => x"7487d302",
  1429 => x"ead9c255",
  1430 => x"9c4c7087",
  1431 => x"c087c702",
  1432 => x"ff05acfb",
  1433 => x"e0c087ed",
  1434 => x"55c1c255",
  1435 => x"d87d97c0",
  1436 => x"a96e4966",
  1437 => x"c887db05",
  1438 => x"66cc4866",
  1439 => x"87ca04a8",
  1440 => x"c14866c8",
  1441 => x"58a6cc80",
  1442 => x"66cc87c8",
  1443 => x"d088c148",
  1444 => x"d8c258a6",
  1445 => x"4c7087ed",
  1446 => x"05acd0c1",
  1447 => x"66d487c8",
  1448 => x"d880c148",
  1449 => x"d0c158a6",
  1450 => x"e6fd02ac",
  1451 => x"a6e0c087",
  1452 => x"7866d848",
  1453 => x"c04866c4",
  1454 => x"05a866e0",
  1455 => x"c087e5c9",
  1456 => x"c048a6e4",
  1457 => x"c080c478",
  1458 => x"c0487478",
  1459 => x"7e7088fb",
  1460 => x"e8c8026e",
  1461 => x"cb486e87",
  1462 => x"6e7e7088",
  1463 => x"87cec102",
  1464 => x"88c9486e",
  1465 => x"026e7e70",
  1466 => x"6e87eac3",
  1467 => x"7088c448",
  1468 => x"ce026e7e",
  1469 => x"c1486e87",
  1470 => x"6e7e7088",
  1471 => x"87d5c302",
  1472 => x"dc87f4c7",
  1473 => x"f0c048a6",
  1474 => x"f6d6c278",
  1475 => x"c04c7087",
  1476 => x"c002acec",
  1477 => x"e0c087c4",
  1478 => x"ecc05ca6",
  1479 => x"cdc002ac",
  1480 => x"ded6c287",
  1481 => x"c04c7087",
  1482 => x"ff05acec",
  1483 => x"ecc087f3",
  1484 => x"c4c002ac",
  1485 => x"cad6c287",
  1486 => x"ca1ec087",
  1487 => x"4966d01e",
  1488 => x"c8c191cb",
  1489 => x"80714866",
  1490 => x"c858a6cc",
  1491 => x"80c44866",
  1492 => x"cc58a6d0",
  1493 => x"ff49bf66",
  1494 => x"c187ebdd",
  1495 => x"d41ede1e",
  1496 => x"ff49bf66",
  1497 => x"d087dfdd",
  1498 => x"c0497086",
  1499 => x"ecc08909",
  1500 => x"e8c059a6",
  1501 => x"a8c04866",
  1502 => x"87eec006",
  1503 => x"4866e8c0",
  1504 => x"c003a8dd",
  1505 => x"66c487e4",
  1506 => x"e8c049bf",
  1507 => x"e0c08166",
  1508 => x"66e8c051",
  1509 => x"c481c149",
  1510 => x"c281bf66",
  1511 => x"e8c051c1",
  1512 => x"81c24966",
  1513 => x"81bf66c4",
  1514 => x"486e51c0",
  1515 => x"78fdcec1",
  1516 => x"81c8496e",
  1517 => x"6e5166d0",
  1518 => x"d481c949",
  1519 => x"496e5166",
  1520 => x"66dc81ca",
  1521 => x"4866d051",
  1522 => x"a6d480c1",
  1523 => x"80d84858",
  1524 => x"e8c478c1",
  1525 => x"deddff87",
  1526 => x"c0497087",
  1527 => x"ff59a6ec",
  1528 => x"7087d4dd",
  1529 => x"a6e0c049",
  1530 => x"4866dc59",
  1531 => x"05a8ecc0",
  1532 => x"dc87cac0",
  1533 => x"e8c048a6",
  1534 => x"c4c07866",
  1535 => x"c2d3c287",
  1536 => x"4966c887",
  1537 => x"c0c191cb",
  1538 => x"80714866",
  1539 => x"4a6e7e70",
  1540 => x"496e82c8",
  1541 => x"e8c081ca",
  1542 => x"66dc5166",
  1543 => x"c081c149",
  1544 => x"c18966e8",
  1545 => x"70307148",
  1546 => x"7189c149",
  1547 => x"d9c47a97",
  1548 => x"c049bfea",
  1549 => x"972966e8",
  1550 => x"71484a6a",
  1551 => x"a6f0c098",
  1552 => x"c4496e58",
  1553 => x"c04d6981",
  1554 => x"c44866e0",
  1555 => x"c002a866",
  1556 => x"a6c487c8",
  1557 => x"c078c048",
  1558 => x"a6c487c5",
  1559 => x"c478c148",
  1560 => x"e0c01e66",
  1561 => x"ff49751e",
  1562 => x"c887dbd9",
  1563 => x"c04c7086",
  1564 => x"c106acb7",
  1565 => x"857487d4",
  1566 => x"7449e0c0",
  1567 => x"c14b7589",
  1568 => x"714ad4e6",
  1569 => x"87e0e0fe",
  1570 => x"e4c085c2",
  1571 => x"80c14866",
  1572 => x"58a6e8c0",
  1573 => x"4966ecc0",
  1574 => x"a97081c1",
  1575 => x"87c8c002",
  1576 => x"c048a6c4",
  1577 => x"87c5c078",
  1578 => x"c148a6c4",
  1579 => x"1e66c478",
  1580 => x"c049a4c2",
  1581 => x"887148e0",
  1582 => x"751e4970",
  1583 => x"c5d8ff49",
  1584 => x"c086c887",
  1585 => x"ff01a8b7",
  1586 => x"e4c087c0",
  1587 => x"d1c00266",
  1588 => x"c9496e87",
  1589 => x"66e4c081",
  1590 => x"c1486e51",
  1591 => x"c078cfd1",
  1592 => x"496e87cc",
  1593 => x"51c281c9",
  1594 => x"d2c1486e",
  1595 => x"e8c078c3",
  1596 => x"78c148a6",
  1597 => x"ff87c6c0",
  1598 => x"7087f6d6",
  1599 => x"66e8c04c",
  1600 => x"87f5c002",
  1601 => x"cc4866c8",
  1602 => x"c004a866",
  1603 => x"66c887cb",
  1604 => x"cc80c148",
  1605 => x"e0c058a6",
  1606 => x"4866cc87",
  1607 => x"a6d088c1",
  1608 => x"87d5c058",
  1609 => x"05acc6c1",
  1610 => x"d087c8c0",
  1611 => x"80c14866",
  1612 => x"ff58a6d4",
  1613 => x"7087fad5",
  1614 => x"4866d44c",
  1615 => x"a6d880c1",
  1616 => x"029c7458",
  1617 => x"c887cbc0",
  1618 => x"c8c14866",
  1619 => x"f204a866",
  1620 => x"d5ff87eb",
  1621 => x"66c887d2",
  1622 => x"03a8c748",
  1623 => x"c487e5c0",
  1624 => x"c048dcd5",
  1625 => x"4966c878",
  1626 => x"c0c191cb",
  1627 => x"a1c48166",
  1628 => x"c04a6a4a",
  1629 => x"66c87952",
  1630 => x"cc80c148",
  1631 => x"a8c758a6",
  1632 => x"87dbff04",
  1633 => x"ff8ed0ff",
  1634 => x"4c87efdf",
  1635 => x"2064616f",
  1636 => x"00202e2a",
  1637 => x"1e00203a",
  1638 => x"4b711e73",
  1639 => x"87c6029b",
  1640 => x"48d8d5c4",
  1641 => x"1ec778c0",
  1642 => x"bfd8d5c4",
  1643 => x"ebc11e49",
  1644 => x"d4c41ee1",
  1645 => x"ed49bfcc",
  1646 => x"86cc87e9",
  1647 => x"bfccd4c4",
  1648 => x"87e3e949",
  1649 => x"c8029b73",
  1650 => x"e1ebc187",
  1651 => x"d8f1c049",
  1652 => x"e9deff87",
  1653 => x"1e731e87",
  1654 => x"4bffc31e",
  1655 => x"fc4ad4ff",
  1656 => x"98c148bf",
  1657 => x"026e7e70",
  1658 => x"ff87fbc0",
  1659 => x"c1c148d0",
  1660 => x"7ad2c278",
  1661 => x"c7c47a73",
  1662 => x"ff4849db",
  1663 => x"73506a80",
  1664 => x"73516a7a",
  1665 => x"6a80c17a",
  1666 => x"6a7a7350",
  1667 => x"6a7a7350",
  1668 => x"6a7a7349",
  1669 => x"6a7a7350",
  1670 => x"e4c7c450",
  1671 => x"d0ff5997",
  1672 => x"78c0c148",
  1673 => x"c7c487d7",
  1674 => x"ff4849db",
  1675 => x"5150c080",
  1676 => x"50c080c1",
  1677 => x"50c150d9",
  1678 => x"c350e2c0",
  1679 => x"e1c7c450",
  1680 => x"f850c048",
  1681 => x"dcff2680",
  1682 => x"cd1e87f4",
  1683 => x"49c187c1",
  1684 => x"fe87c4fd",
  1685 => x"7087ebe3",
  1686 => x"87cd0298",
  1687 => x"87e6ecfe",
  1688 => x"c4029870",
  1689 => x"c24ac187",
  1690 => x"724ac087",
  1691 => x"87ce059a",
  1692 => x"eac11ec0",
  1693 => x"fbc049df",
  1694 => x"86c487d6",
  1695 => x"edc187fe",
  1696 => x"1ec087e8",
  1697 => x"49eaeac1",
  1698 => x"87c4fbc0",
  1699 => x"d0c21ec0",
  1700 => x"497087cf",
  1701 => x"87f8fac0",
  1702 => x"f887ffc2",
  1703 => x"534f268e",
  1704 => x"61662044",
  1705 => x"64656c69",
  1706 => x"6f42002e",
  1707 => x"6e69746f",
  1708 => x"2e2e2e67",
  1709 => x"d5c41e00",
  1710 => x"78c048d8",
  1711 => x"48ccd4c4",
  1712 => x"c5fe78c0",
  1713 => x"c7d2c287",
  1714 => x"2648c087",
  1715 => x"0100004f",
  1716 => x"80000000",
  1717 => x"69784520",
  1718 => x"20800074",
  1719 => x"6b636142",
  1720 => x"0013ff00",
  1721 => x"00456c00",
  1722 => x"00000000",
  1723 => x"000013ff",
  1724 => x"0000458a",
  1725 => x"ff000000",
  1726 => x"a8000013",
  1727 => x"00000045",
  1728 => x"13ff0000",
  1729 => x"45c60000",
  1730 => x"00000000",
  1731 => x"0013ff00",
  1732 => x"0045e400",
  1733 => x"00000000",
  1734 => x"000013ff",
  1735 => x"00004602",
  1736 => x"ff000000",
  1737 => x"20000013",
  1738 => x"00000046",
  1739 => x"13ff0000",
  1740 => x"00000000",
  1741 => x"00000000",
  1742 => x"00149400",
  1743 => x"00000000",
  1744 => x"00000000",
  1745 => x"48f0fe1e",
  1746 => x"09cd78c0",
  1747 => x"4f260979",
  1748 => x"f0fe1e1e",
  1749 => x"26487ebf",
  1750 => x"fe1e4f26",
  1751 => x"78c148f0",
  1752 => x"fe1e4f26",
  1753 => x"78c048f0",
  1754 => x"711e4f26",
  1755 => x"7a97c04a",
  1756 => x"c049a2c1",
  1757 => x"49a2ca51",
  1758 => x"a2cb51c0",
  1759 => x"2651c049",
  1760 => x"5b5e0e4f",
  1761 => x"86f00e5c",
  1762 => x"a4ca4c71",
  1763 => x"7e699749",
  1764 => x"974ba4cb",
  1765 => x"a6c8486b",
  1766 => x"cc80c158",
  1767 => x"98c758a6",
  1768 => x"6e58a6d0",
  1769 => x"a866cc48",
  1770 => x"9787db05",
  1771 => x"6b977e69",
  1772 => x"58a6c848",
  1773 => x"a6cc80c1",
  1774 => x"d098c758",
  1775 => x"486e58a6",
  1776 => x"02a866cc",
  1777 => x"d9fe87e5",
  1778 => x"4aa4cc87",
  1779 => x"72496b97",
  1780 => x"66dc49a1",
  1781 => x"7e6b9751",
  1782 => x"80c1486e",
  1783 => x"c758a6c8",
  1784 => x"58a6cc98",
  1785 => x"c37b9770",
  1786 => x"edfd87d2",
  1787 => x"c28ef087",
  1788 => x"264d2687",
  1789 => x"264b264c",
  1790 => x"5b5e0e4f",
  1791 => x"f40e5d5c",
  1792 => x"974d7186",
  1793 => x"a5c17e6d",
  1794 => x"486c974c",
  1795 => x"6e58a6c8",
  1796 => x"a866c448",
  1797 => x"ff87c505",
  1798 => x"87e6c048",
  1799 => x"c287c3fd",
  1800 => x"6c9749a5",
  1801 => x"4ba3714b",
  1802 => x"974b6b97",
  1803 => x"486e7e6c",
  1804 => x"a6c880c1",
  1805 => x"cc98c758",
  1806 => x"977058a6",
  1807 => x"87dafc7c",
  1808 => x"8ef44873",
  1809 => x"0e87eafe",
  1810 => x"0e5c5b5e",
  1811 => x"4c7186f4",
  1812 => x"c34a66d8",
  1813 => x"a4c29aff",
  1814 => x"496c974b",
  1815 => x"7249a173",
  1816 => x"7e6c9751",
  1817 => x"80c1486e",
  1818 => x"c758a6c8",
  1819 => x"58a6cc98",
  1820 => x"8ef45470",
  1821 => x"1e87fcfd",
  1822 => x"699786f0",
  1823 => x"4aa1c17e",
  1824 => x"c8486a97",
  1825 => x"486e58a6",
  1826 => x"a8b766c4",
  1827 => x"9787d304",
  1828 => x"6a977e69",
  1829 => x"58a6c848",
  1830 => x"66c4486e",
  1831 => x"58a6cc88",
  1832 => x"7e1187d6",
  1833 => x"80c8486e",
  1834 => x"481258a6",
  1835 => x"c458a6cc",
  1836 => x"66c84866",
  1837 => x"58a6d088",
  1838 => x"4f268ef0",
  1839 => x"f41e731e",
  1840 => x"87defa86",
  1841 => x"494bbfe0",
  1842 => x"99c0e0c0",
  1843 => x"7387cb02",
  1844 => x"fed8c41e",
  1845 => x"87effd49",
  1846 => x"497386c4",
  1847 => x"0299c0d0",
  1848 => x"c487c0c1",
  1849 => x"bf97c8d9",
  1850 => x"c9d9c47e",
  1851 => x"c848bf97",
  1852 => x"486e58a6",
  1853 => x"02a866c4",
  1854 => x"c487e8c0",
  1855 => x"bf97c8d9",
  1856 => x"cad9c449",
  1857 => x"e0481181",
  1858 => x"d9c47808",
  1859 => x"7ebf97c8",
  1860 => x"80c1486e",
  1861 => x"c758a6c8",
  1862 => x"58a6cc98",
  1863 => x"48c8d9c4",
  1864 => x"e45066c8",
  1865 => x"c0494bbf",
  1866 => x"0299c0e0",
  1867 => x"1e7387cb",
  1868 => x"49d2d9c4",
  1869 => x"c487d0fc",
  1870 => x"d0497386",
  1871 => x"c10299c0",
  1872 => x"d9c487c0",
  1873 => x"7ebf97dc",
  1874 => x"97ddd9c4",
  1875 => x"a6c848bf",
  1876 => x"c4486e58",
  1877 => x"c002a866",
  1878 => x"d9c487e8",
  1879 => x"49bf97dc",
  1880 => x"81ded9c4",
  1881 => x"08e44811",
  1882 => x"dcd9c478",
  1883 => x"6e7ebf97",
  1884 => x"c880c148",
  1885 => x"98c758a6",
  1886 => x"c458a6cc",
  1887 => x"c848dcd9",
  1888 => x"cbf75066",
  1889 => x"f77e7087",
  1890 => x"8ef487d0",
  1891 => x"1e87e6f9",
  1892 => x"49fed8c4",
  1893 => x"c487d3f7",
  1894 => x"f749d2d9",
  1895 => x"f2c187cc",
  1896 => x"dff649fc",
  1897 => x"87d0c387",
  1898 => x"5e0e4f26",
  1899 => x"710e5c5b",
  1900 => x"fed8c44c",
  1901 => x"87c1f949",
  1902 => x"b7c04a70",
  1903 => x"e3c204aa",
  1904 => x"aaf0c387",
  1905 => x"c187c905",
  1906 => x"c148f0f9",
  1907 => x"87c4c278",
  1908 => x"05aae0c3",
  1909 => x"f9c187c9",
  1910 => x"78c148f4",
  1911 => x"c187f5c1",
  1912 => x"02bff4f9",
  1913 => x"c0c287c6",
  1914 => x"87c24ba2",
  1915 => x"9c744b72",
  1916 => x"c187d205",
  1917 => x"1ebff0f9",
  1918 => x"bff4f9c1",
  1919 => x"c149721e",
  1920 => x"c887d1f8",
  1921 => x"f0f9c186",
  1922 => x"e0c002bf",
  1923 => x"c4497387",
  1924 => x"c19129b7",
  1925 => x"7381c7fb",
  1926 => x"c29acf4a",
  1927 => x"7248c192",
  1928 => x"ff4a7030",
  1929 => x"694872ba",
  1930 => x"db797098",
  1931 => x"c4497387",
  1932 => x"c19129b7",
  1933 => x"7381c7fb",
  1934 => x"c29acf4a",
  1935 => x"7248c392",
  1936 => x"484a7030",
  1937 => x"7970b069",
  1938 => x"48f4f9c1",
  1939 => x"f9c178c0",
  1940 => x"78c048f0",
  1941 => x"49fed8c4",
  1942 => x"7087def6",
  1943 => x"aab7c04a",
  1944 => x"87ddfd03",
  1945 => x"87c248c0",
  1946 => x"4c264d26",
  1947 => x"4f264b26",
  1948 => x"00000000",
  1949 => x"00000000",
  1950 => x"724ac01e",
  1951 => x"c191c449",
  1952 => x"c081c7fb",
  1953 => x"d082c179",
  1954 => x"ee04aab7",
  1955 => x"0e4f2687",
  1956 => x"5d5c5b5e",
  1957 => x"f34d710e",
  1958 => x"4a7587c8",
  1959 => x"922ab7c4",
  1960 => x"82c7fbc1",
  1961 => x"9ccf4c75",
  1962 => x"496a94c2",
  1963 => x"c32b744b",
  1964 => x"7448c29b",
  1965 => x"ff4c7030",
  1966 => x"714874bc",
  1967 => x"f27a7098",
  1968 => x"487387d8",
  1969 => x"0087e1fe",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00000000",
  1984 => x"00000000",
  1985 => x"0e000000",
  1986 => x"5d5c5b5e",
  1987 => x"9a4a710e",
  1988 => x"c287c602",
  1989 => x"c048e8c2",
  1990 => x"e8c2c278",
  1991 => x"c6c105bf",
  1992 => x"d2d9c487",
  1993 => x"87d1f349",
  1994 => x"04a8b7c0",
  1995 => x"d9c487cd",
  1996 => x"c4f349d2",
  1997 => x"a8b7c087",
  1998 => x"c287f303",
  1999 => x"49bfe8c2",
  2000 => x"48e8c2c2",
  2001 => x"c278a1c1",
  2002 => x"1181f8c2",
  2003 => x"f0c2c248",
  2004 => x"f0c2c258",
  2005 => x"c078c048",
  2006 => x"e9c049f2",
  2007 => x"497087cf",
  2008 => x"59ead9c4",
  2009 => x"c287f9c4",
  2010 => x"02bff0c2",
  2011 => x"c487f2c1",
  2012 => x"f249d2d9",
  2013 => x"b7c087c3",
  2014 => x"87cd04a8",
  2015 => x"bff0c2c2",
  2016 => x"c288c148",
  2017 => x"db58f4c2",
  2018 => x"e6d9c487",
  2019 => x"e8c049bf",
  2020 => x"987087e7",
  2021 => x"c487cd02",
  2022 => x"ef49d2d9",
  2023 => x"c2c287cc",
  2024 => x"78c048e8",
  2025 => x"bfecc2c2",
  2026 => x"87f4c305",
  2027 => x"bff0c2c2",
  2028 => x"87ecc305",
  2029 => x"bfe8c2c2",
  2030 => x"e8c2c249",
  2031 => x"78a1c148",
  2032 => x"81f8c2c2",
  2033 => x"c2494b11",
  2034 => x"c00299c0",
  2035 => x"487387cc",
  2036 => x"c298ffc1",
  2037 => x"c358f4c2",
  2038 => x"c2c287c6",
  2039 => x"ffc25bf0",
  2040 => x"ecc2c287",
  2041 => x"dbc102bf",
  2042 => x"e6d9c487",
  2043 => x"e7c049bf",
  2044 => x"987087c7",
  2045 => x"87e8c202",
  2046 => x"bfe8c2c2",
  2047 => x"e8c2c249",
  2048 => x"78a1c148",
  2049 => x"81f8c2c2",
  2050 => x"1e496997",
  2051 => x"49d2d9c4",
  2052 => x"c487eeed",
  2053 => x"ecc2c286",
  2054 => x"89c149bf",
  2055 => x"59f0c2c2",
  2056 => x"48f0c2c2",
  2057 => x"997178c1",
  2058 => x"87c6c002",
  2059 => x"c04cf2c0",
  2060 => x"dcd787c3",
  2061 => x"c049744c",
  2062 => x"7087f2e5",
  2063 => x"ead9c449",
  2064 => x"87dcc159",
  2065 => x"49d2d9c4",
  2066 => x"7087ecf0",
  2067 => x"c0029b4b",
  2068 => x"c2c287ee",
  2069 => x"abb7bff4",
  2070 => x"87e4c003",
  2071 => x"bfe6d9c4",
  2072 => x"d4e5c049",
  2073 => x"02987087",
  2074 => x"c787f5c0",
  2075 => x"f4c2c248",
  2076 => x"c2c288bf",
  2077 => x"d9c458f8",
  2078 => x"edeb49d2",
  2079 => x"87e0c087",
  2080 => x"c049dcd7",
  2081 => x"7087e6e4",
  2082 => x"ead9c449",
  2083 => x"f4c2c259",
  2084 => x"abb74abf",
  2085 => x"87c8c004",
  2086 => x"d5f1c149",
  2087 => x"87e4fe87",
  2088 => x"4c264d26",
  2089 => x"4f264b26",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000004",
  2094 => x"0882ff01",
  2095 => x"64f3c8f3",
  2096 => x"01f250f3",
  2097 => x"00f40181",
  2098 => x"48d0ff1e",
  2099 => x"7178e1c8",
  2100 => x"08d4ff48",
  2101 => x"1e4f2678",
  2102 => x"c848d0ff",
  2103 => x"487178e1",
  2104 => x"7808d4ff",
  2105 => x"ff4866c4",
  2106 => x"267808d4",
  2107 => x"4a711e4f",
  2108 => x"1e4966c4",
  2109 => x"deff4972",
  2110 => x"48d0ff87",
  2111 => x"2678e0c0",
  2112 => x"731e4f26",
  2113 => x"c84b711e",
  2114 => x"731e4966",
  2115 => x"a2e0c14a",
  2116 => x"87d9ff49",
  2117 => x"2687c426",
  2118 => x"264c264d",
  2119 => x"1e4f264b",
  2120 => x"4b711e73",
  2121 => x"fe49e2c0",
  2122 => x"4ac787de",
  2123 => x"d4ff4813",
  2124 => x"49727808",
  2125 => x"99718ac1",
  2126 => x"ff87f105",
  2127 => x"e0c048d0",
  2128 => x"87d7ff78",
  2129 => x"5c5b5e0e",
  2130 => x"4c710e5d",
  2131 => x"bfead9c4",
  2132 => x"2b744b4d",
  2133 => x"c19b66d0",
  2134 => x"ab66d483",
  2135 => x"c087c204",
  2136 => x"d04a744b",
  2137 => x"31724966",
  2138 => x"9975b9ff",
  2139 => x"30724873",
  2140 => x"71484a70",
  2141 => x"eed9c4b0",
  2142 => x"efecc158",
  2143 => x"264d2687",
  2144 => x"264b264c",
  2145 => x"d0ff1e4f",
  2146 => x"78c9c848",
  2147 => x"d4ff4871",
  2148 => x"4f267808",
  2149 => x"494a711e",
  2150 => x"d0ff87eb",
  2151 => x"2678c848",
  2152 => x"1e731e4f",
  2153 => x"d9c44b71",
  2154 => x"c302bffa",
  2155 => x"87ebc287",
  2156 => x"c848d0ff",
  2157 => x"497378c9",
  2158 => x"ffb1e0c0",
  2159 => x"787148d4",
  2160 => x"48eed9c4",
  2161 => x"66c878c0",
  2162 => x"c387c502",
  2163 => x"87c249ff",
  2164 => x"d9c449c0",
  2165 => x"66cc59f6",
  2166 => x"c587c602",
  2167 => x"c44ad5d5",
  2168 => x"ffffcf87",
  2169 => x"fad9c44a",
  2170 => x"fad9c45a",
  2171 => x"c478c148",
  2172 => x"264d2687",
  2173 => x"264b264c",
  2174 => x"5b5e0e4f",
  2175 => x"710e5d5c",
  2176 => x"f6d9c44a",
  2177 => x"9a724cbf",
  2178 => x"4987cb02",
  2179 => x"c6c291c8",
  2180 => x"83714bd7",
  2181 => x"cac287c4",
  2182 => x"4dc04bd7",
  2183 => x"99744913",
  2184 => x"bff2d9c4",
  2185 => x"48d4ffb9",
  2186 => x"b7c17871",
  2187 => x"b7c8852c",
  2188 => x"87e804ad",
  2189 => x"bfeed9c4",
  2190 => x"c480c848",
  2191 => x"fe58f2d9",
  2192 => x"731e87ef",
  2193 => x"134b711e",
  2194 => x"cb029a4a",
  2195 => x"fe497287",
  2196 => x"4a1387e7",
  2197 => x"87f5059a",
  2198 => x"1e87dafe",
  2199 => x"bfeed9c4",
  2200 => x"eed9c449",
  2201 => x"78a1c148",
  2202 => x"a9b7c0c4",
  2203 => x"ff87db03",
  2204 => x"d9c448d4",
  2205 => x"c478bff2",
  2206 => x"49bfeed9",
  2207 => x"48eed9c4",
  2208 => x"c478a1c1",
  2209 => x"04a9b7c0",
  2210 => x"d0ff87e5",
  2211 => x"c478c848",
  2212 => x"c048fad9",
  2213 => x"004f2678",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"5f5f0000",
  2217 => x"00000000",
  2218 => x"03000303",
  2219 => x"14000003",
  2220 => x"7f147f7f",
  2221 => x"0000147f",
  2222 => x"6b6b2e24",
  2223 => x"4c00123a",
  2224 => x"6c18366a",
  2225 => x"30003256",
  2226 => x"77594f7e",
  2227 => x"0040683a",
  2228 => x"03070400",
  2229 => x"00000000",
  2230 => x"633e1c00",
  2231 => x"00000041",
  2232 => x"3e634100",
  2233 => x"0800001c",
  2234 => x"1c1c3e2a",
  2235 => x"00082a3e",
  2236 => x"3e3e0808",
  2237 => x"00000808",
  2238 => x"60e08000",
  2239 => x"00000000",
  2240 => x"08080808",
  2241 => x"00000808",
  2242 => x"60600000",
  2243 => x"40000000",
  2244 => x"0c183060",
  2245 => x"00010306",
  2246 => x"4d597f3e",
  2247 => x"00003e7f",
  2248 => x"7f7f0604",
  2249 => x"00000000",
  2250 => x"59716342",
  2251 => x"0000464f",
  2252 => x"49496322",
  2253 => x"1800367f",
  2254 => x"7f13161c",
  2255 => x"0000107f",
  2256 => x"45456727",
  2257 => x"0000397d",
  2258 => x"494b7e3c",
  2259 => x"00003079",
  2260 => x"79710101",
  2261 => x"0000070f",
  2262 => x"49497f36",
  2263 => x"0000367f",
  2264 => x"69494f06",
  2265 => x"00001e3f",
  2266 => x"66660000",
  2267 => x"00000000",
  2268 => x"66e68000",
  2269 => x"00000000",
  2270 => x"14140808",
  2271 => x"00002222",
  2272 => x"14141414",
  2273 => x"00001414",
  2274 => x"14142222",
  2275 => x"00000808",
  2276 => x"59510302",
  2277 => x"3e00060f",
  2278 => x"555d417f",
  2279 => x"00001e1f",
  2280 => x"09097f7e",
  2281 => x"00007e7f",
  2282 => x"49497f7f",
  2283 => x"0000367f",
  2284 => x"41633e1c",
  2285 => x"00004141",
  2286 => x"63417f7f",
  2287 => x"00001c3e",
  2288 => x"49497f7f",
  2289 => x"00004141",
  2290 => x"09097f7f",
  2291 => x"00000101",
  2292 => x"49417f3e",
  2293 => x"00007a7b",
  2294 => x"08087f7f",
  2295 => x"00007f7f",
  2296 => x"7f7f4100",
  2297 => x"00000041",
  2298 => x"40406020",
  2299 => x"7f003f7f",
  2300 => x"361c087f",
  2301 => x"00004163",
  2302 => x"40407f7f",
  2303 => x"7f004040",
  2304 => x"060c067f",
  2305 => x"7f007f7f",
  2306 => x"180c067f",
  2307 => x"00007f7f",
  2308 => x"41417f3e",
  2309 => x"00003e7f",
  2310 => x"09097f7f",
  2311 => x"3e00060f",
  2312 => x"7f61417f",
  2313 => x"0000407e",
  2314 => x"19097f7f",
  2315 => x"0000667f",
  2316 => x"594d6f26",
  2317 => x"0000327b",
  2318 => x"7f7f0101",
  2319 => x"00000101",
  2320 => x"40407f3f",
  2321 => x"00003f7f",
  2322 => x"70703f0f",
  2323 => x"7f000f3f",
  2324 => x"3018307f",
  2325 => x"41007f7f",
  2326 => x"1c1c3663",
  2327 => x"01416336",
  2328 => x"7c7c0603",
  2329 => x"61010306",
  2330 => x"474d5971",
  2331 => x"00004143",
  2332 => x"417f7f00",
  2333 => x"01000041",
  2334 => x"180c0603",
  2335 => x"00406030",
  2336 => x"7f414100",
  2337 => x"0800007f",
  2338 => x"0603060c",
  2339 => x"8000080c",
  2340 => x"80808080",
  2341 => x"00008080",
  2342 => x"07030000",
  2343 => x"00000004",
  2344 => x"54547420",
  2345 => x"0000787c",
  2346 => x"44447f7f",
  2347 => x"0000387c",
  2348 => x"44447c38",
  2349 => x"00000044",
  2350 => x"44447c38",
  2351 => x"00007f7f",
  2352 => x"54547c38",
  2353 => x"0000185c",
  2354 => x"057f7e04",
  2355 => x"00000005",
  2356 => x"a4a4bc18",
  2357 => x"00007cfc",
  2358 => x"04047f7f",
  2359 => x"0000787c",
  2360 => x"7d3d0000",
  2361 => x"00000040",
  2362 => x"fd808080",
  2363 => x"0000007d",
  2364 => x"38107f7f",
  2365 => x"0000446c",
  2366 => x"7f3f0000",
  2367 => x"7c000040",
  2368 => x"0c180c7c",
  2369 => x"0000787c",
  2370 => x"04047c7c",
  2371 => x"0000787c",
  2372 => x"44447c38",
  2373 => x"0000387c",
  2374 => x"2424fcfc",
  2375 => x"0000183c",
  2376 => x"24243c18",
  2377 => x"0000fcfc",
  2378 => x"04047c7c",
  2379 => x"0000080c",
  2380 => x"54545c48",
  2381 => x"00002074",
  2382 => x"447f3f04",
  2383 => x"00000044",
  2384 => x"40407c3c",
  2385 => x"00007c7c",
  2386 => x"60603c1c",
  2387 => x"3c001c3c",
  2388 => x"6030607c",
  2389 => x"44003c7c",
  2390 => x"3810386c",
  2391 => x"0000446c",
  2392 => x"60e0bc1c",
  2393 => x"00001c3c",
  2394 => x"5c746444",
  2395 => x"0000444c",
  2396 => x"773e0808",
  2397 => x"00004141",
  2398 => x"7f7f0000",
  2399 => x"00000000",
  2400 => x"3e774141",
  2401 => x"02000808",
  2402 => x"02030101",
  2403 => x"7f000102",
  2404 => x"7f7f7f7f",
  2405 => x"08007f7f",
  2406 => x"3e1c1c08",
  2407 => x"7f7f7f3e",
  2408 => x"1c3e3e7f",
  2409 => x"0008081c",
  2410 => x"7c7c1810",
  2411 => x"00001018",
  2412 => x"7c7c3010",
  2413 => x"10001030",
  2414 => x"78606030",
  2415 => x"4200061e",
  2416 => x"3c183c66",
  2417 => x"78004266",
  2418 => x"c6c26a38",
  2419 => x"6000386c",
  2420 => x"00600000",
  2421 => x"0e006000",
  2422 => x"5d5c5b5e",
  2423 => x"4c711e0e",
  2424 => x"bfcbdac4",
  2425 => x"c04bc04d",
  2426 => x"02ab741e",
  2427 => x"a6c487c7",
  2428 => x"c578c048",
  2429 => x"48a6c487",
  2430 => x"66c478c1",
  2431 => x"ee49731e",
  2432 => x"86c887df",
  2433 => x"ef49e0c0",
  2434 => x"a5c487ef",
  2435 => x"f0496a4a",
  2436 => x"c6f187f0",
  2437 => x"c185cb87",
  2438 => x"abb7c883",
  2439 => x"87c7ff04",
  2440 => x"264d2626",
  2441 => x"264b264c",
  2442 => x"4a711e4f",
  2443 => x"5acfdac4",
  2444 => x"48cfdac4",
  2445 => x"fe4978c7",
  2446 => x"4f2687dd",
  2447 => x"711e731e",
  2448 => x"aab7c04a",
  2449 => x"c287d303",
  2450 => x"05bfe5e6",
  2451 => x"4bc187c4",
  2452 => x"4bc087c2",
  2453 => x"5be9e6c2",
  2454 => x"e6c287c4",
  2455 => x"e6c25ae9",
  2456 => x"c14abfe5",
  2457 => x"a2c0c19a",
  2458 => x"87e8ec49",
  2459 => x"e6c248fc",
  2460 => x"fe78bfe5",
  2461 => x"c21e87ef",
  2462 => x"48bfe5e6",
  2463 => x"711e4f26",
  2464 => x"1e66c44a",
  2465 => x"f9e94972",
  2466 => x"4f262687",
  2467 => x"e5e6c21e",
  2468 => x"d8c149bf",
  2469 => x"dac487c5",
  2470 => x"bfe848c3",
  2471 => x"ffd9c478",
  2472 => x"78bfec48",
  2473 => x"bfc3dac4",
  2474 => x"ffc3494a",
  2475 => x"2ab7c899",
  2476 => x"b0714872",
  2477 => x"58cbdac4",
  2478 => x"5e0e4f26",
  2479 => x"0e5d5c5b",
  2480 => x"c7ff4b71",
  2481 => x"fed9c487",
  2482 => x"7350c048",
  2483 => x"fedeff49",
  2484 => x"4c497087",
  2485 => x"eecb9cc2",
  2486 => x"87d1cb49",
  2487 => x"c44d4970",
  2488 => x"bf97fed9",
  2489 => x"87e4c105",
  2490 => x"c44966d0",
  2491 => x"99bfc7da",
  2492 => x"d487d705",
  2493 => x"d9c44966",
  2494 => x"0599bfff",
  2495 => x"497387cc",
  2496 => x"87cbdeff",
  2497 => x"c1029870",
  2498 => x"4cc187c2",
  2499 => x"7587fdfd",
  2500 => x"87e5ca49",
  2501 => x"c6029870",
  2502 => x"fed9c487",
  2503 => x"c450c148",
  2504 => x"bf97fed9",
  2505 => x"87e4c005",
  2506 => x"bfc7dac4",
  2507 => x"9966d049",
  2508 => x"87d6ff05",
  2509 => x"bfffd9c4",
  2510 => x"9966d449",
  2511 => x"87caff05",
  2512 => x"ddff4973",
  2513 => x"987087c9",
  2514 => x"87fefe05",
  2515 => x"d0fb4874",
  2516 => x"5b5e0e87",
  2517 => x"f40e5d5c",
  2518 => x"4c4dc086",
  2519 => x"c47ebfec",
  2520 => x"dac448a6",
  2521 => x"c178bfcb",
  2522 => x"c31ec01e",
  2523 => x"c9fd49fc",
  2524 => x"7086c887",
  2525 => x"87ce0298",
  2526 => x"fffa49ff",
  2527 => x"49dac187",
  2528 => x"87cbdcff",
  2529 => x"d9c44dc1",
  2530 => x"02bf97fe",
  2531 => x"f8c087c4",
  2532 => x"dac487ef",
  2533 => x"c24bbfc3",
  2534 => x"05bfe5e6",
  2535 => x"c387ebc0",
  2536 => x"dbff49fd",
  2537 => x"fac387e9",
  2538 => x"e2dbff49",
  2539 => x"c3497387",
  2540 => x"1e7199ff",
  2541 => x"c5fb49c0",
  2542 => x"c8497387",
  2543 => x"1e7129b7",
  2544 => x"f9fa49c1",
  2545 => x"c686c887",
  2546 => x"dac487c1",
  2547 => x"9b4bbfc7",
  2548 => x"c287dd02",
  2549 => x"49bfe1e6",
  2550 => x"7087dec7",
  2551 => x"87c40598",
  2552 => x"87d24bc0",
  2553 => x"c749e0c2",
  2554 => x"e6c287c3",
  2555 => x"87c658e5",
  2556 => x"48e1e6c2",
  2557 => x"497378c0",
  2558 => x"ce0599c2",
  2559 => x"49ebc387",
  2560 => x"87cbdaff",
  2561 => x"99c24970",
  2562 => x"fb87c202",
  2563 => x"c149734c",
  2564 => x"87ce0599",
  2565 => x"ff49f4c3",
  2566 => x"7087f4d9",
  2567 => x"0299c249",
  2568 => x"4cfa87c2",
  2569 => x"99c84973",
  2570 => x"c387ce05",
  2571 => x"d9ff49f5",
  2572 => x"497087dd",
  2573 => x"d50299c2",
  2574 => x"cfdac487",
  2575 => x"87ca02bf",
  2576 => x"c488c148",
  2577 => x"c058d3da",
  2578 => x"4cff87c2",
  2579 => x"49734dc1",
  2580 => x"ce0599c4",
  2581 => x"49f2c387",
  2582 => x"87f3d8ff",
  2583 => x"99c24970",
  2584 => x"c487dc02",
  2585 => x"7ebfcfda",
  2586 => x"a8b7c748",
  2587 => x"87cbc003",
  2588 => x"80c1486e",
  2589 => x"58d3dac4",
  2590 => x"fe87c2c0",
  2591 => x"c34dc14c",
  2592 => x"d8ff49fd",
  2593 => x"497087c9",
  2594 => x"c00299c2",
  2595 => x"dac487d5",
  2596 => x"c002bfcf",
  2597 => x"dac487c9",
  2598 => x"78c048cf",
  2599 => x"fd87c2c0",
  2600 => x"c34dc14c",
  2601 => x"d7ff49fa",
  2602 => x"497087e5",
  2603 => x"c00299c2",
  2604 => x"dac487d9",
  2605 => x"c748bfcf",
  2606 => x"c003a8b7",
  2607 => x"dac487c9",
  2608 => x"78c748cf",
  2609 => x"fc87c2c0",
  2610 => x"c04dc14c",
  2611 => x"c003acb7",
  2612 => x"66c487d1",
  2613 => x"82d8c14a",
  2614 => x"c6c0026a",
  2615 => x"744b6a87",
  2616 => x"c00f7349",
  2617 => x"1ef0c31e",
  2618 => x"f749dac1",
  2619 => x"86c887cc",
  2620 => x"c0029870",
  2621 => x"a6c887e2",
  2622 => x"cfdac448",
  2623 => x"66c878bf",
  2624 => x"c491cb49",
  2625 => x"80714866",
  2626 => x"bf6e7e70",
  2627 => x"87c8c002",
  2628 => x"c84bbf6e",
  2629 => x"0f734966",
  2630 => x"c0029d75",
  2631 => x"dac487c8",
  2632 => x"f249bfcf",
  2633 => x"e6c287f1",
  2634 => x"c002bfe9",
  2635 => x"c24987dd",
  2636 => x"987087c7",
  2637 => x"87d3c002",
  2638 => x"bfcfdac4",
  2639 => x"87d7f249",
  2640 => x"f7f349c0",
  2641 => x"e9e6c287",
  2642 => x"f478c048",
  2643 => x"87d1f38e",
  2644 => x"5c5b5e0e",
  2645 => x"711e0e5d",
  2646 => x"cbdac44c",
  2647 => x"cdc149bf",
  2648 => x"d1c14da1",
  2649 => x"747e6981",
  2650 => x"87cf029c",
  2651 => x"744ba5c4",
  2652 => x"cbdac47b",
  2653 => x"f0f249bf",
  2654 => x"747b6e87",
  2655 => x"87c4059c",
  2656 => x"87c24bc0",
  2657 => x"49734bc1",
  2658 => x"d487f1f2",
  2659 => x"87c70266",
  2660 => x"7087da49",
  2661 => x"c087c24a",
  2662 => x"ede6c24a",
  2663 => x"c0f2265a",
  2664 => x"00000087",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"4a711e00",
  2668 => x"49bfc8ff",
  2669 => x"2648a172",
  2670 => x"c8ff1e4f",
  2671 => x"c0fe89bf",
  2672 => x"c0c0c0c0",
  2673 => x"87c401a9",
  2674 => x"87c24ac0",
  2675 => x"48724ac1",
  2676 => x"5e0e4f26",
  2677 => x"0e5d5c5b",
  2678 => x"d4ff4b71",
  2679 => x"4866d04c",
  2680 => x"49d678c0",
  2681 => x"87e0dbff",
  2682 => x"6c7cffc3",
  2683 => x"99ffc349",
  2684 => x"c3494d71",
  2685 => x"e0c199f0",
  2686 => x"87cb05a9",
  2687 => x"6c7cffc3",
  2688 => x"d098c348",
  2689 => x"c3780866",
  2690 => x"4a6c7cff",
  2691 => x"c331c849",
  2692 => x"4a6c7cff",
  2693 => x"4972b271",
  2694 => x"ffc331c8",
  2695 => x"714a6c7c",
  2696 => x"c84972b2",
  2697 => x"7cffc331",
  2698 => x"b2714a6c",
  2699 => x"c048d0ff",
  2700 => x"9b7378e0",
  2701 => x"7287c202",
  2702 => x"2648757b",
  2703 => x"264c264d",
  2704 => x"1e4f264b",
  2705 => x"5e0e4f26",
  2706 => x"f80e5c5b",
  2707 => x"c81e7686",
  2708 => x"fdfd49a6",
  2709 => x"7086c487",
  2710 => x"c2486e4b",
  2711 => x"f4c203a8",
  2712 => x"c34a7387",
  2713 => x"d0c19af0",
  2714 => x"87c702aa",
  2715 => x"05aae0c1",
  2716 => x"7387e2c2",
  2717 => x"0299c849",
  2718 => x"c6ff87c3",
  2719 => x"c34c7387",
  2720 => x"05acc29c",
  2721 => x"c487c4c1",
  2722 => x"31c94966",
  2723 => x"66c41e71",
  2724 => x"92c8c14a",
  2725 => x"49d3dac4",
  2726 => x"c2fe8172",
  2727 => x"49d887d6",
  2728 => x"87e4d8ff",
  2729 => x"c41ec0c8",
  2730 => x"fd49dac7",
  2731 => x"ff87e2da",
  2732 => x"e0c048d0",
  2733 => x"dac7c478",
  2734 => x"4a66cc1e",
  2735 => x"c492c8c1",
  2736 => x"7249d3da",
  2737 => x"e0fdfd81",
  2738 => x"c186cc87",
  2739 => x"c4c105ac",
  2740 => x"4966c487",
  2741 => x"1e7131c9",
  2742 => x"c14a66c4",
  2743 => x"dac492c8",
  2744 => x"817249d3",
  2745 => x"87ccc1fe",
  2746 => x"1edac7c4",
  2747 => x"c14a66c8",
  2748 => x"dac492c8",
  2749 => x"817249d3",
  2750 => x"87defbfd",
  2751 => x"d7ff49d7",
  2752 => x"c0c887c6",
  2753 => x"dac7c41e",
  2754 => x"ddd8fd49",
  2755 => x"ff86cc87",
  2756 => x"e0c048d0",
  2757 => x"fc8ef878",
  2758 => x"5e0e87e3",
  2759 => x"0e5d5c5b",
  2760 => x"ff4d711e",
  2761 => x"66d44cd4",
  2762 => x"b7c3487e",
  2763 => x"87c506a8",
  2764 => x"e3c148c0",
  2765 => x"fe497587",
  2766 => x"7587e6d0",
  2767 => x"4b66c41e",
  2768 => x"c493c8c1",
  2769 => x"7383d3da",
  2770 => x"e6f4fd49",
  2771 => x"6b83c887",
  2772 => x"48d0ff4b",
  2773 => x"dd78e1c8",
  2774 => x"c349737c",
  2775 => x"7c7199ff",
  2776 => x"b7c84973",
  2777 => x"99ffc329",
  2778 => x"49737c71",
  2779 => x"c329b7d0",
  2780 => x"7c7199ff",
  2781 => x"b7d84973",
  2782 => x"c07c7129",
  2783 => x"7c7c7c7c",
  2784 => x"7c7c7c7c",
  2785 => x"7c7c7c7c",
  2786 => x"c478e0c0",
  2787 => x"49dc1e66",
  2788 => x"87d9d5ff",
  2789 => x"487386c8",
  2790 => x"87dffa26",
  2791 => x"4ad4ff1e",
  2792 => x"c848d0ff",
  2793 => x"f0c378c5",
  2794 => x"c07a717a",
  2795 => x"7a7a7a7a",
  2796 => x"4f2678c4",
  2797 => x"4ad4ff1e",
  2798 => x"c848d0ff",
  2799 => x"7ac078c5",
  2800 => x"7ac0496a",
  2801 => x"7a7a7a7a",
  2802 => x"487178c4",
  2803 => x"731e4f26",
  2804 => x"c84b711e",
  2805 => x"87db0266",
  2806 => x"c14a6b97",
  2807 => x"699749a3",
  2808 => x"51727b97",
  2809 => x"c24866c8",
  2810 => x"58a6cc88",
  2811 => x"987083c2",
  2812 => x"c487e505",
  2813 => x"264d2687",
  2814 => x"264b264c",
  2815 => x"5b5e0e4f",
  2816 => x"e80e5d5c",
  2817 => x"59a6cc86",
  2818 => x"4d66e8c0",
  2819 => x"c495dcc1",
  2820 => x"c185e3dc",
  2821 => x"c47ea5c8",
  2822 => x"ccc148a6",
  2823 => x"66c478a5",
  2824 => x"bf6e4cbf",
  2825 => x"85d0c194",
  2826 => x"66c8946d",
  2827 => x"c84ac04b",
  2828 => x"d2fd49c0",
  2829 => x"66c887c2",
  2830 => x"9fc0c148",
  2831 => x"4966c878",
  2832 => x"bf6e81c2",
  2833 => x"66c8799f",
  2834 => x"c481c649",
  2835 => x"799fbf66",
  2836 => x"cc4966c8",
  2837 => x"799f6d81",
  2838 => x"d44866c8",
  2839 => x"58a6d080",
  2840 => x"48e9f4c2",
  2841 => x"d44966cc",
  2842 => x"41204aa1",
  2843 => x"f905aa71",
  2844 => x"4866c887",
  2845 => x"d480eec0",
  2846 => x"f4c258a6",
  2847 => x"66d048fe",
  2848 => x"4aa1c849",
  2849 => x"aa714120",
  2850 => x"c887f905",
  2851 => x"f6c04866",
  2852 => x"58a6d880",
  2853 => x"48c7f5c2",
  2854 => x"c04966d4",
  2855 => x"204aa1e8",
  2856 => x"05aa7141",
  2857 => x"e8c087f9",
  2858 => x"4966d81e",
  2859 => x"cc87dffc",
  2860 => x"dec14966",
  2861 => x"d0c0c881",
  2862 => x"66cc799f",
  2863 => x"81e2c149",
  2864 => x"799fc0c8",
  2865 => x"c14966cc",
  2866 => x"9fc181ea",
  2867 => x"4966cc79",
  2868 => x"c481ecc1",
  2869 => x"799fbf66",
  2870 => x"c14966cc",
  2871 => x"66c881ee",
  2872 => x"cc799fbf",
  2873 => x"f0c14966",
  2874 => x"799f6d81",
  2875 => x"ffcf4b74",
  2876 => x"4a739bff",
  2877 => x"c14966cc",
  2878 => x"9f7281f2",
  2879 => x"d04a7479",
  2880 => x"ffffcf2a",
  2881 => x"cc4c729a",
  2882 => x"f4c14966",
  2883 => x"799f7481",
  2884 => x"4966cc73",
  2885 => x"7381f8c1",
  2886 => x"cc72799f",
  2887 => x"fac14966",
  2888 => x"799f7281",
  2889 => x"ccfb8ee4",
  2890 => x"544d6987",
  2891 => x"694d6953",
  2892 => x"484d696e",
  2893 => x"66617267",
  2894 => x"20696c64",
  2895 => x"312e0065",
  2896 => x"20203030",
  2897 => x"59002020",
  2898 => x"42555141",
  2899 => x"20202045",
  2900 => x"20202020",
  2901 => x"20202020",
  2902 => x"20202020",
  2903 => x"20202020",
  2904 => x"20202020",
  2905 => x"20202020",
  2906 => x"20202020",
  2907 => x"00202020",
  2908 => x"711e731e",
  2909 => x"0266d44b",
  2910 => x"66c887d4",
  2911 => x"7331d849",
  2912 => x"7232c84a",
  2913 => x"66cc49a1",
  2914 => x"c0487181",
  2915 => x"66d087e3",
  2916 => x"91dcc149",
  2917 => x"81e3dcc4",
  2918 => x"4aa1ccc1",
  2919 => x"92734a6a",
  2920 => x"c18266c8",
  2921 => x"496981d0",
  2922 => x"66cc9172",
  2923 => x"7189c181",
  2924 => x"87c5f948",
  2925 => x"ff4a711e",
  2926 => x"d0ff49d4",
  2927 => x"78c5c848",
  2928 => x"c079d0c2",
  2929 => x"79797979",
  2930 => x"79797979",
  2931 => x"79c07972",
  2932 => x"c07966c4",
  2933 => x"7966c879",
  2934 => x"66cc79c0",
  2935 => x"d079c079",
  2936 => x"79c07966",
  2937 => x"c47966d4",
  2938 => x"1e4f2678",
  2939 => x"a2c64a71",
  2940 => x"49699749",
  2941 => x"7199f0c3",
  2942 => x"1e1ec01e",
  2943 => x"1ec01ec1",
  2944 => x"87f0fe49",
  2945 => x"f649d0c2",
  2946 => x"8eec87d2",
  2947 => x"c01e4f26",
  2948 => x"1e1e1e1e",
  2949 => x"fe49c11e",
  2950 => x"d0c287da",
  2951 => x"87fcf549",
  2952 => x"4f268eec",
  2953 => x"ff4a711e",
  2954 => x"c5c848d0",
  2955 => x"48d4ff78",
  2956 => x"c078e0c2",
  2957 => x"78787878",
  2958 => x"1ec0c878",
  2959 => x"cbfd4972",
  2960 => x"d0ff87e8",
  2961 => x"2678c448",
  2962 => x"5e0e4f26",
  2963 => x"0e5d5c5b",
  2964 => x"4a7186f8",
  2965 => x"c14ba2c2",
  2966 => x"a2c37b97",
  2967 => x"7c97c14c",
  2968 => x"51c049a2",
  2969 => x"c04da2c4",
  2970 => x"a2c57d97",
  2971 => x"c0486e7e",
  2972 => x"48a6c450",
  2973 => x"c478a2c6",
  2974 => x"50c04866",
  2975 => x"c41e66d8",
  2976 => x"f549dac7",
  2977 => x"66c887f7",
  2978 => x"1e49bf97",
  2979 => x"bf9766c8",
  2980 => x"49151e49",
  2981 => x"1e49141e",
  2982 => x"c01e4913",
  2983 => x"87d4fc49",
  2984 => x"f7f349c8",
  2985 => x"dac7c487",
  2986 => x"87f8fd49",
  2987 => x"f349d0c2",
  2988 => x"8ee087ea",
  2989 => x"1e87fef4",
  2990 => x"a2c64a71",
  2991 => x"49699749",
  2992 => x"49a2c51e",
  2993 => x"1e496997",
  2994 => x"9749a2c4",
  2995 => x"c31e4969",
  2996 => x"699749a2",
  2997 => x"a2c21e49",
  2998 => x"49699749",
  2999 => x"fb49c01e",
  3000 => x"d0c287d2",
  3001 => x"87f4f249",
  3002 => x"4f268eec",
  3003 => x"711e731e",
  3004 => x"4aa3c24b",
  3005 => x"c14966c8",
  3006 => x"dcc491dc",
  3007 => x"d4c181e3",
  3008 => x"c2791281",
  3009 => x"d3f249d0",
  3010 => x"87edf387",
  3011 => x"711e731e",
  3012 => x"49a3c64b",
  3013 => x"1e496997",
  3014 => x"9749a3c5",
  3015 => x"c41e4969",
  3016 => x"699749a3",
  3017 => x"a3c31e49",
  3018 => x"49699749",
  3019 => x"49a3c21e",
  3020 => x"1e496997",
  3021 => x"124aa3c1",
  3022 => x"87f8f949",
  3023 => x"f149d0c2",
  3024 => x"8eec87da",
  3025 => x"0e87f2f2",
  3026 => x"5d5c5b5e",
  3027 => x"7e711e0e",
  3028 => x"81c2496e",
  3029 => x"6e7997c1",
  3030 => x"c183c34b",
  3031 => x"4a6e7b97",
  3032 => x"97c082c1",
  3033 => x"c44c6e7a",
  3034 => x"7c97c084",
  3035 => x"85c54d6e",
  3036 => x"4d6e55c0",
  3037 => x"6d9785c6",
  3038 => x"1ec01e4d",
  3039 => x"1e4c6c97",
  3040 => x"1e4b6b97",
  3041 => x"1e496997",
  3042 => x"e7f84912",
  3043 => x"49d0c287",
  3044 => x"e887c9f0",
  3045 => x"87ddf18e",
  3046 => x"5c5b5e0e",
  3047 => x"dcff0e5d",
  3048 => x"c34b7186",
  3049 => x"4c1149a3",
  3050 => x"c54aa3c4",
  3051 => x"699749a3",
  3052 => x"9731c849",
  3053 => x"71484a6a",
  3054 => x"58a6d4b0",
  3055 => x"6e7ea3c6",
  3056 => x"4d49bf97",
  3057 => x"48719dcf",
  3058 => x"d898c0c1",
  3059 => x"f04858a6",
  3060 => x"78a3c280",
  3061 => x"bf9766c4",
  3062 => x"58a6d048",
  3063 => x"c01e66d4",
  3064 => x"741e66f8",
  3065 => x"c01e751e",
  3066 => x"f64966e0",
  3067 => x"86d087c2",
  3068 => x"a6dc4970",
  3069 => x"0266cc59",
  3070 => x"c087e4c5",
  3071 => x"c50266f8",
  3072 => x"4a66cc87",
  3073 => x"4ac187c2",
  3074 => x"f8c04b72",
  3075 => x"87db0266",
  3076 => x"4966f4c0",
  3077 => x"c491dcc1",
  3078 => x"c181e3dc",
  3079 => x"a6c881d4",
  3080 => x"c8786948",
  3081 => x"06aab766",
  3082 => x"c84b87c1",
  3083 => x"87eced49",
  3084 => x"7087c1ee",
  3085 => x"0599c449",
  3086 => x"f7ed87ca",
  3087 => x"c4497087",
  3088 => x"87f60299",
  3089 => x"88c14873",
  3090 => x"58a6e0c0",
  3091 => x"dc80ec48",
  3092 => x"9b737866",
  3093 => x"87d0c102",
  3094 => x"c14866cc",
  3095 => x"f0c002a8",
  3096 => x"66f4c087",
  3097 => x"91dcc149",
  3098 => x"4ae3dcc4",
  3099 => x"d0c18271",
  3100 => x"ac6949a2",
  3101 => x"c187d805",
  3102 => x"ccc1854c",
  3103 => x"ad6949a2",
  3104 => x"c087ce05",
  3105 => x"4866d04d",
  3106 => x"a6d480c1",
  3107 => x"c187c258",
  3108 => x"4866cc84",
  3109 => x"a6d088c1",
  3110 => x"4966c858",
  3111 => x"cc88c148",
  3112 => x"997158a6",
  3113 => x"87f0fe05",
  3114 => x"d90266d4",
  3115 => x"d8497387",
  3116 => x"4a718166",
  3117 => x"729affc3",
  3118 => x"c84a714c",
  3119 => x"a6d42ab7",
  3120 => x"29b7d85a",
  3121 => x"976e4d71",
  3122 => x"f0c349bf",
  3123 => x"71b17599",
  3124 => x"4966d41e",
  3125 => x"7129b7c8",
  3126 => x"1e66d81e",
  3127 => x"66d41e74",
  3128 => x"1e49bf97",
  3129 => x"cbf349c0",
  3130 => x"d086d487",
  3131 => x"87ecea49",
  3132 => x"4966f4c0",
  3133 => x"c491dcc1",
  3134 => x"7148e3dc",
  3135 => x"58a6cc80",
  3136 => x"c84966c8",
  3137 => x"c1026981",
  3138 => x"e0c087ca",
  3139 => x"66dc48a6",
  3140 => x"029b7378",
  3141 => x"d887c2c1",
  3142 => x"31c94966",
  3143 => x"66cc1e71",
  3144 => x"cfe8fd49",
  3145 => x"d01ec087",
  3146 => x"e2fd4966",
  3147 => x"1ec187ec",
  3148 => x"fd4966d4",
  3149 => x"cc87c9e1",
  3150 => x"4866d886",
  3151 => x"a6dc80c1",
  3152 => x"66e0c058",
  3153 => x"88c14849",
  3154 => x"58a6e4c0",
  3155 => x"ff059971",
  3156 => x"87c587c5",
  3157 => x"c3e949c9",
  3158 => x"0566cc87",
  3159 => x"c287dcfa",
  3160 => x"f7e849c0",
  3161 => x"8edcff87",
  3162 => x"0e87caea",
  3163 => x"5d5c5b5e",
  3164 => x"7186e00e",
  3165 => x"49a4c34c",
  3166 => x"a6d44811",
  3167 => x"4aa4c458",
  3168 => x"9749a4c5",
  3169 => x"31c84969",
  3170 => x"484a6a97",
  3171 => x"a6d8b071",
  3172 => x"7ea4c658",
  3173 => x"49bf976e",
  3174 => x"719dcf4d",
  3175 => x"98c0c148",
  3176 => x"4858a6dc",
  3177 => x"a4c280ec",
  3178 => x"9766c478",
  3179 => x"66d84bbf",
  3180 => x"66f4c01e",
  3181 => x"1e66d81e",
  3182 => x"e4c01e75",
  3183 => x"efee4966",
  3184 => x"7086d087",
  3185 => x"a6e0c049",
  3186 => x"059b7359",
  3187 => x"c0c487c3",
  3188 => x"e749c44b",
  3189 => x"66dc87c6",
  3190 => x"7131c949",
  3191 => x"66f4c01e",
  3192 => x"91dcc149",
  3193 => x"48e3dcc4",
  3194 => x"a6d48071",
  3195 => x"4966d058",
  3196 => x"87c0e5fd",
  3197 => x"9b7386c4",
  3198 => x"87dfc402",
  3199 => x"0266f4c0",
  3200 => x"4a7387c4",
  3201 => x"4ac187c2",
  3202 => x"f4c04c72",
  3203 => x"87d30266",
  3204 => x"c14966cc",
  3205 => x"a6c881d4",
  3206 => x"c8786948",
  3207 => x"06aab766",
  3208 => x"744c87c1",
  3209 => x"d5c2029c",
  3210 => x"87c8e687",
  3211 => x"99c84970",
  3212 => x"e587ca05",
  3213 => x"497087fe",
  3214 => x"f60299c8",
  3215 => x"48d0ff87",
  3216 => x"ff78c5c8",
  3217 => x"f0c248d4",
  3218 => x"7878c078",
  3219 => x"c8787878",
  3220 => x"c7c41ec0",
  3221 => x"fbfc49da",
  3222 => x"d0ff87f7",
  3223 => x"c478c448",
  3224 => x"d41edac7",
  3225 => x"defd4966",
  3226 => x"1ec187ff",
  3227 => x"fd4966d8",
  3228 => x"cc87cddc",
  3229 => x"4866dc86",
  3230 => x"e0c080c1",
  3231 => x"abc158a6",
  3232 => x"87f3c002",
  3233 => x"c14966cc",
  3234 => x"66d081d0",
  3235 => x"05a86948",
  3236 => x"a6d087dd",
  3237 => x"8578c148",
  3238 => x"c14966cc",
  3239 => x"ad6981cc",
  3240 => x"c087d405",
  3241 => x"4866d44d",
  3242 => x"a6d880c1",
  3243 => x"d087c858",
  3244 => x"80c14866",
  3245 => x"c158a6d4",
  3246 => x"fd058c8b",
  3247 => x"66d887eb",
  3248 => x"dc87da02",
  3249 => x"ffc34966",
  3250 => x"59a6d499",
  3251 => x"c84966dc",
  3252 => x"a6d829b7",
  3253 => x"4966dc59",
  3254 => x"7129b7d8",
  3255 => x"bf976e4d",
  3256 => x"99f0c349",
  3257 => x"1e71b175",
  3258 => x"c84966d8",
  3259 => x"1e7129b7",
  3260 => x"dc1e66dc",
  3261 => x"66d41e66",
  3262 => x"1e49bf97",
  3263 => x"f3ea49c0",
  3264 => x"7386d487",
  3265 => x"87c7029b",
  3266 => x"cfe249d0",
  3267 => x"c287c687",
  3268 => x"c7e249d0",
  3269 => x"059b7387",
  3270 => x"e087e1fb",
  3271 => x"87d5e38e",
  3272 => x"5c5b5e0e",
  3273 => x"86e40e5d",
  3274 => x"a6cc4a71",
  3275 => x"78ffc048",
  3276 => x"ffc180c4",
  3277 => x"c380c478",
  3278 => x"80c478ff",
  3279 => x"a2c878c0",
  3280 => x"c9496949",
  3281 => x"9d4d7129",
  3282 => x"87eec202",
  3283 => x"a6cc4cc0",
  3284 => x"c2026b4b",
  3285 => x"497487ca",
  3286 => x"a17391c4",
  3287 => x"c87e6949",
  3288 => x"78c448a6",
  3289 => x"6e4966c8",
  3290 => x"721e7191",
  3291 => x"4a09751e",
  3292 => x"87c5f6fc",
  3293 => x"49264a26",
  3294 => x"c458a6c8",
  3295 => x"b7c0c0c0",
  3296 => x"87cb01ad",
  3297 => x"a8b7ffcf",
  3298 => x"87fdc006",
  3299 => x"c487ebc0",
  3300 => x"ffc34866",
  3301 => x"04a8b7ff",
  3302 => x"c487eec0",
  3303 => x"ffc74866",
  3304 => x"03a8b7ff",
  3305 => x"66c887c9",
  3306 => x"a8b7c548",
  3307 => x"c487da03",
  3308 => x"ffcf4866",
  3309 => x"06a8b7ff",
  3310 => x"66c887cf",
  3311 => x"cc80c148",
  3312 => x"b7d058a6",
  3313 => x"dbfe06a8",
  3314 => x"4866c887",
  3315 => x"06a8b7d0",
  3316 => x"84c187ce",
  3317 => x"91c44974",
  3318 => x"6949a173",
  3319 => x"87f6fd05",
  3320 => x"49a2c8c1",
  3321 => x"c17966c4",
  3322 => x"c849a2cc",
  3323 => x"d0c17966",
  3324 => x"796e49a2",
  3325 => x"49a2d4c1",
  3326 => x"8ee479c1",
  3327 => x"87f5dfff",
  3328 => x"c449c01e",
  3329 => x"02bfebdc",
  3330 => x"49c187c2",
  3331 => x"bfc7dec4",
  3332 => x"c287c202",
  3333 => x"48d0ffb1",
  3334 => x"ff78c5c8",
  3335 => x"fac348d4",
  3336 => x"ff787178",
  3337 => x"78c448d0",
  3338 => x"731e4f26",
  3339 => x"1e4a711e",
  3340 => x"c14966cc",
  3341 => x"dcc491dc",
  3342 => x"83714be3",
  3343 => x"d0fd4973",
  3344 => x"86c487f1",
  3345 => x"c5029870",
  3346 => x"fb497387",
  3347 => x"effe87d2",
  3348 => x"e4deff87",
  3349 => x"5b5e0e87",
  3350 => x"f40e5d5c",
  3351 => x"d3ddff86",
  3352 => x"c4497087",
  3353 => x"d2c50299",
  3354 => x"48d0ff87",
  3355 => x"ff78c5c8",
  3356 => x"c0c248d4",
  3357 => x"7878c078",
  3358 => x"4d787878",
  3359 => x"c048d4ff",
  3360 => x"a54a7678",
  3361 => x"bfd4ff49",
  3362 => x"d4ff7997",
  3363 => x"6878c048",
  3364 => x"c885c151",
  3365 => x"e304adb7",
  3366 => x"48d0ff87",
  3367 => x"97c678c4",
  3368 => x"a6cc4866",
  3369 => x"d04c7058",
  3370 => x"2cb7c49c",
  3371 => x"dcc14974",
  3372 => x"e3dcc491",
  3373 => x"6981c881",
  3374 => x"c287ca05",
  3375 => x"dbff49d1",
  3376 => x"f6c387da",
  3377 => x"6697c787",
  3378 => x"f0c3494b",
  3379 => x"05a9d099",
  3380 => x"1e7487cc",
  3381 => x"d2e44972",
  3382 => x"c386c487",
  3383 => x"d0c287dd",
  3384 => x"87c805ab",
  3385 => x"e5e44972",
  3386 => x"87cfc387",
  3387 => x"05abecc3",
  3388 => x"1ec087ce",
  3389 => x"49721e74",
  3390 => x"c887cfe5",
  3391 => x"87fbc286",
  3392 => x"05abd1c2",
  3393 => x"1e7487cc",
  3394 => x"eae64972",
  3395 => x"c286c487",
  3396 => x"c6c387e9",
  3397 => x"87cc05ab",
  3398 => x"49721e74",
  3399 => x"c487cde7",
  3400 => x"87d7c286",
  3401 => x"05abe0c0",
  3402 => x"1ec087ce",
  3403 => x"49721e74",
  3404 => x"c887e5e9",
  3405 => x"87c3c286",
  3406 => x"05abc4c3",
  3407 => x"1ec187ce",
  3408 => x"49721e74",
  3409 => x"c887d1e9",
  3410 => x"87efc186",
  3411 => x"05abf0c0",
  3412 => x"1ec087ce",
  3413 => x"49721e74",
  3414 => x"c887d0f0",
  3415 => x"87dbc186",
  3416 => x"05abc5c3",
  3417 => x"1ec187ce",
  3418 => x"49721e74",
  3419 => x"c887fcef",
  3420 => x"87c7c186",
  3421 => x"cc05abc8",
  3422 => x"721e7487",
  3423 => x"87c7e749",
  3424 => x"f6c086c4",
  3425 => x"059b7387",
  3426 => x"1e7487cc",
  3427 => x"fbe54972",
  3428 => x"c086c487",
  3429 => x"66c887e5",
  3430 => x"6697c91e",
  3431 => x"97cc1e49",
  3432 => x"cf1e4966",
  3433 => x"1e496697",
  3434 => x"496697d2",
  3435 => x"e049c41e",
  3436 => x"86d487c2",
  3437 => x"ff49d1c2",
  3438 => x"f487e1d7",
  3439 => x"f4d8ff8e",
  3440 => x"d8c31e87",
  3441 => x"c149bfcf",
  3442 => x"d3d8c3b9",
  3443 => x"48d4ff59",
  3444 => x"ff78ffc3",
  3445 => x"e1c048d0",
  3446 => x"48d4ff78",
  3447 => x"31c478c1",
  3448 => x"d0ff7871",
  3449 => x"78e0c048",
  3450 => x"c31e4f26",
  3451 => x"c41ec3d8",
  3452 => x"fd49d0d4",
  3453 => x"c487fcc9",
  3454 => x"02987086",
  3455 => x"c0ff87c3",
  3456 => x"314f2687",
  3457 => x"5a484b35",
  3458 => x"43202020",
  3459 => x"00004746",
  3460 => x"1e000000",
  3461 => x"87dec1ff",
  3462 => x"87c6d5fe",
  3463 => x"c24966c4",
  3464 => x"cd0299c0",
  3465 => x"1ee0c387",
  3466 => x"49fed8c4",
  3467 => x"87d7d8fe",
  3468 => x"66c486c4",
  3469 => x"99c0c449",
  3470 => x"c387cd02",
  3471 => x"d8c41ef0",
  3472 => x"d8fe49fe",
  3473 => x"86c487c1",
  3474 => x"c14966c4",
  3475 => x"1e7199ff",
  3476 => x"49fed8c4",
  3477 => x"87efd7fe",
  3478 => x"87fed3fe",
  3479 => x"0e4f2626",
  3480 => x"5d5c5b5e",
  3481 => x"86d8ff0e",
  3482 => x"dfc47ec0",
  3483 => x"c249bfdf",
  3484 => x"721e7181",
  3485 => x"fc4ac61e",
  3486 => x"7187fee9",
  3487 => x"264a2648",
  3488 => x"58a6c849",
  3489 => x"bfdfdfc4",
  3490 => x"7181c449",
  3491 => x"c61e721e",
  3492 => x"e4e9fc4a",
  3493 => x"26487187",
  3494 => x"cc49264a",
  3495 => x"e4c358a6",
  3496 => x"ff49bff2",
  3497 => x"7087d2cc",
  3498 => x"fac90298",
  3499 => x"49e0c087",
  3500 => x"87f9cbff",
  3501 => x"e4c34970",
  3502 => x"4cc059f6",
  3503 => x"91c44974",
  3504 => x"6981d0fe",
  3505 => x"c449744a",
  3506 => x"81bfdfdf",
  3507 => x"dfc491c4",
  3508 => x"797281eb",
  3509 => x"87d2029a",
  3510 => x"89c14972",
  3511 => x"486e9a71",
  3512 => x"7e7080c1",
  3513 => x"ff059a72",
  3514 => x"84c187ee",
  3515 => x"04acb7c2",
  3516 => x"6e87c9ff",
  3517 => x"b7fcc048",
  3518 => x"eac804a8",
  3519 => x"744cc087",
  3520 => x"8266c44a",
  3521 => x"dfc492c4",
  3522 => x"497482eb",
  3523 => x"c48166c8",
  3524 => x"ebdfc491",
  3525 => x"694a6a81",
  3526 => x"74b97249",
  3527 => x"dfdfc44b",
  3528 => x"93c483bf",
  3529 => x"83ebdfc4",
  3530 => x"4872ba6b",
  3531 => x"a6d49871",
  3532 => x"c4497458",
  3533 => x"81bfdfdf",
  3534 => x"dfc491c4",
  3535 => x"7e6981eb",
  3536 => x"c048a6d4",
  3537 => x"5ca6d078",
  3538 => x"d04cffc3",
  3539 => x"29df4966",
  3540 => x"87e2c602",
  3541 => x"c04a66cc",
  3542 => x"66d492e0",
  3543 => x"48ffc082",
  3544 => x"4a708872",
  3545 => x"c048a6d8",
  3546 => x"c080c478",
  3547 => x"df496e78",
  3548 => x"a6e4c029",
  3549 => x"dbdfc459",
  3550 => x"7278c148",
  3551 => x"b731c349",
  3552 => x"c0b1722a",
  3553 => x"91c499ff",
  3554 => x"4dc8c0c4",
  3555 => x"4b6d8571",
  3556 => x"c0c0c449",
  3557 => x"87d70299",
  3558 => x"0266e0c0",
  3559 => x"c887c7c0",
  3560 => x"c578c080",
  3561 => x"dfc487d0",
  3562 => x"78c148e3",
  3563 => x"c087c7c5",
  3564 => x"d80266e0",
  3565 => x"c2497387",
  3566 => x"0299c0c0",
  3567 => x"d087c3c0",
  3568 => x"486d2bb7",
  3569 => x"98fffffd",
  3570 => x"fac07d70",
  3571 => x"e3dfc487",
  3572 => x"f2c002bf",
  3573 => x"d0487387",
  3574 => x"e8c028b7",
  3575 => x"987058a6",
  3576 => x"87e3c002",
  3577 => x"bfe7dfc4",
  3578 => x"c0e0c049",
  3579 => x"cac00299",
  3580 => x"c0497087",
  3581 => x"0299c0e0",
  3582 => x"6d87ccc0",
  3583 => x"c0c0c248",
  3584 => x"c07d70b0",
  3585 => x"734b66e4",
  3586 => x"c0c0c849",
  3587 => x"c5c20299",
  3588 => x"e7dfc487",
  3589 => x"c0cc4abf",
  3590 => x"cfc0029a",
  3591 => x"8ac0c487",
  3592 => x"87d7c002",
  3593 => x"f8c0028a",
  3594 => x"87dcc187",
  3595 => x"99744973",
  3596 => x"ffc391c2",
  3597 => x"4b1181fc",
  3598 => x"7387dbc1",
  3599 => x"c2997449",
  3600 => x"fcffc391",
  3601 => x"1181c181",
  3602 => x"66e0c04b",
  3603 => x"87c8c002",
  3604 => x"d248a6dc",
  3605 => x"87fec078",
  3606 => x"c448a6d8",
  3607 => x"f5c078d2",
  3608 => x"74497387",
  3609 => x"c391c299",
  3610 => x"c181fcff",
  3611 => x"c04b1181",
  3612 => x"c00266e0",
  3613 => x"a6dc87c9",
  3614 => x"78d9c148",
  3615 => x"d887d7c0",
  3616 => x"d9c548a6",
  3617 => x"87cec078",
  3618 => x"99744973",
  3619 => x"ffc391c2",
  3620 => x"81c181fc",
  3621 => x"e0c04b11",
  3622 => x"dbc00266",
  3623 => x"ff497387",
  3624 => x"c0fcc7b9",
  3625 => x"c4487199",
  3626 => x"98bfe7df",
  3627 => x"58ebdfc4",
  3628 => x"c0c49b74",
  3629 => x"87d3c0b3",
  3630 => x"fcc74973",
  3631 => x"487199c0",
  3632 => x"bfe7dfc4",
  3633 => x"ebdfc4b0",
  3634 => x"d89b7458",
  3635 => x"cac00266",
  3636 => x"dfc41e87",
  3637 => x"faf449db",
  3638 => x"7386c487",
  3639 => x"dbdfc41e",
  3640 => x"87eff449",
  3641 => x"66dc86c4",
  3642 => x"87cac002",
  3643 => x"dbdfc41e",
  3644 => x"87dff449",
  3645 => x"66d086c4",
  3646 => x"d430c148",
  3647 => x"486e58a6",
  3648 => x"7e7030c1",
  3649 => x"c14866d4",
  3650 => x"58a6d880",
  3651 => x"a8b7e0c0",
  3652 => x"87f7f804",
  3653 => x"c14c66cc",
  3654 => x"acb7c284",
  3655 => x"87dff704",
  3656 => x"48dfdfc4",
  3657 => x"ff7866c4",
  3658 => x"4d268ed8",
  3659 => x"4b264c26",
  3660 => x"00004f26",
  3661 => x"c01e0000",
  3662 => x"c449724a",
  3663 => x"ebdfc491",
  3664 => x"c179ff81",
  3665 => x"aab7c682",
  3666 => x"c487ee04",
  3667 => x"c048dfdf",
  3668 => x"26784040",
  3669 => x"711e1e4f",
  3670 => x"c7e0c44a",
  3671 => x"c1487ebf",
  3672 => x"cbe0c480",
  3673 => x"81c44958",
  3674 => x"5172816e",
  3675 => x"e0c498cf",
  3676 => x"dc4858cb",
  3677 => x"c840c680",
  3678 => x"66cc7866",
  3679 => x"ecc0ff49",
  3680 => x"c4497087",
  3681 => x"2659e3e0",
  3682 => x"731e4f26",
  3683 => x"494a711e",
  3684 => x"c00299c1",
  3685 => x"66c887eb",
  3686 => x"0299c149",
  3687 => x"c0c387c5",
  3688 => x"c387c34b",
  3689 => x"c8c34bd0",
  3690 => x"731ec41e",
  3691 => x"feb1c749",
  3692 => x"c8c387e3",
  3693 => x"dc1ec41e",
  3694 => x"b1734966",
  3695 => x"d087d6fe",
  3696 => x"87eafd86",
  3697 => x"5c5b5e0e",
  3698 => x"86f80e5d",
  3699 => x"bfdfe0c4",
  3700 => x"e4fffe49",
  3701 => x"7e497087",
  3702 => x"dbfe49c4",
  3703 => x"d4ff87ea",
  3704 => x"78ffc348",
  3705 => x"ffc34968",
  3706 => x"48a6c478",
  3707 => x"78bfd4ff",
  3708 => x"c048d0ff",
  3709 => x"e1c278e0",
  3710 => x"f1c205a9",
  3711 => x"4a66c487",
  3712 => x"028ae0c0",
  3713 => x"d087c3c2",
  3714 => x"d3c2028a",
  3715 => x"028ac187",
  3716 => x"8a87cdc2",
  3717 => x"87c8c202",
  3718 => x"c3c2028a",
  3719 => x"028acc87",
  3720 => x"c287f5c1",
  3721 => x"c0028afe",
  3722 => x"8ac187fd",
  3723 => x"8a87d502",
  3724 => x"87fac105",
  3725 => x"c11ec8c3",
  3726 => x"49ffc31e",
  3727 => x"c887d6fc",
  3728 => x"87eac186",
  3729 => x"bfe3e0c4",
  3730 => x"05a8c148",
  3731 => x"c8c387d0",
  3732 => x"c31ec21e",
  3733 => x"fcfb49fe",
  3734 => x"c186c887",
  3735 => x"e0c487d0",
  3736 => x"78c048e3",
  3737 => x"c487c7c1",
  3738 => x"48bfe3e0",
  3739 => x"d005a8c2",
  3740 => x"1ec8c387",
  3741 => x"fdc31ec3",
  3742 => x"87d9fb49",
  3743 => x"edc086c8",
  3744 => x"e3e0c487",
  3745 => x"c078c048",
  3746 => x"1ec087e4",
  3747 => x"c1c21ec3",
  3748 => x"87c1fb49",
  3749 => x"87d686c8",
  3750 => x"48e3e0c4",
  3751 => x"87ce78c3",
  3752 => x"c34866c4",
  3753 => x"dfe0c498",
  3754 => x"80c84858",
  3755 => x"e0c478c3",
  3756 => x"c24bbfe3",
  3757 => x"e4c0028b",
  3758 => x"028bc187",
  3759 => x"8b87f3c0",
  3760 => x"8b87cc02",
  3761 => x"8b87c802",
  3762 => x"87eac302",
  3763 => x"6e87e5c4",
  3764 => x"87e0c402",
  3765 => x"48e3e0c4",
  3766 => x"d7c478c3",
  3767 => x"c4026e87",
  3768 => x"c8c387d2",
  3769 => x"c31ec11e",
  3770 => x"e8f949ff",
  3771 => x"c486c887",
  3772 => x"e0c487c2",
  3773 => x"c249bfdb",
  3774 => x"f3c10299",
  3775 => x"ebe0c487",
  3776 => x"c8c005bf",
  3777 => x"efe0c487",
  3778 => x"e3c102bf",
  3779 => x"ebe0c487",
  3780 => x"ff4c4dbf",
  3781 => x"03adb7c0",
  3782 => x"4c87c1c0",
  3783 => x"acb7ffc0",
  3784 => x"87c1c006",
  3785 => x"7448754c",
  3786 => x"efe0c488",
  3787 => x"1ec8c358",
  3788 => x"49741ec4",
  3789 => x"f899ffc1",
  3790 => x"86c887db",
  3791 => x"bfefe0c4",
  3792 => x"8c0cc04c",
  3793 => x"acb7c0ff",
  3794 => x"87c1c003",
  3795 => x"b7ffc04c",
  3796 => x"c1c006ac",
  3797 => x"e0c44c87",
  3798 => x"7448bfef",
  3799 => x"f3e0c480",
  3800 => x"1ec8c358",
  3801 => x"49741ec5",
  3802 => x"f799ffc1",
  3803 => x"86c887e7",
  3804 => x"bfdbe0c4",
  3805 => x"0299c149",
  3806 => x"c487fbc0",
  3807 => x"4cbff3e0",
  3808 => x"bfd0f0c3",
  3809 => x"c0bb744b",
  3810 => x"731e741e",
  3811 => x"87faf749",
  3812 => x"b72bb7c1",
  3813 => x"741ec22c",
  3814 => x"f749731e",
  3815 => x"b7c187ec",
  3816 => x"1e2cb72b",
  3817 => x"49731e74",
  3818 => x"d887dff7",
  3819 => x"d0f0c386",
  3820 => x"f3e0c448",
  3821 => x"e0c478bf",
  3822 => x"c448bfc7",
  3823 => x"a8bfc3e0",
  3824 => x"87f0c002",
  3825 => x"80c1487e",
  3826 => x"58c7e0c4",
  3827 => x"6e83c84b",
  3828 => x"4b6b9783",
  3829 => x"e0c498cf",
  3830 => x"49c558c7",
  3831 => x"87e8d3fe",
  3832 => x"7348d4ff",
  3833 => x"48d0ff78",
  3834 => x"c478e0c0",
  3835 => x"c448e3e0",
  3836 => x"78bfe7e0",
  3837 => x"bfc7e0c4",
  3838 => x"c3e0c448",
  3839 => x"c005a8bf",
  3840 => x"7ec087c5",
  3841 => x"c187c2c0",
  3842 => x"f8486e7e",
  3843 => x"87daf48e",
  3844 => x"00000000",
  3845 => x"5c5b5e0e",
  3846 => x"4b710e5d",
  3847 => x"e0c44cc0",
  3848 => x"c405bfdb",
  3849 => x"c24dc187",
  3850 => x"754dc087",
  3851 => x"0599c149",
  3852 => x"d087e5c1",
  3853 => x"87c30266",
  3854 => x"73b3c0c2",
  3855 => x"cec9fe49",
  3856 => x"d44a7087",
  3857 => x"87c60566",
  3858 => x"c1059a72",
  3859 => x"fec387ca",
  3860 => x"817449d3",
  3861 => x"029a4a11",
  3862 => x"7387fdc0",
  3863 => x"f2c005aa",
  3864 => x"0266d487",
  3865 => x"d0c387c5",
  3866 => x"c387c34d",
  3867 => x"c8c34dc0",
  3868 => x"741ec41e",
  3869 => x"2ab7c44a",
  3870 => x"b1754972",
  3871 => x"c387d6f3",
  3872 => x"1ec41ec8",
  3873 => x"9acf4a74",
  3874 => x"b1754972",
  3875 => x"d087c6f3",
  3876 => x"c187c586",
  3877 => x"87f6fe84",
  3878 => x"1e87cff2",
  3879 => x"4b711e73",
  3880 => x"7387fce6",
  3881 => x"c1c4fe49",
  3882 => x"87c2f287",
  3883 => x"fe49c11e",
  3884 => x"ff87d5d0",
  3885 => x"d9c448d4",
  3886 => x"ff78bfea",
  3887 => x"e0c048d0",
  3888 => x"1e4f2678",
  3889 => x"e0c44ac0",
  3890 => x"ca02bff7",
  3891 => x"e0c44987",
  3892 => x"a1c148f7",
  3893 => x"724a1178",
  3894 => x"87c6059a",
  3895 => x"48f7e0c4",
  3896 => x"487278c0",
  3897 => x"c41e4f26",
  3898 => x"c448f7e0",
  3899 => x"78bfc8c4",
  3900 => x"5e0e4f26",
  3901 => x"0e5d5c5b",
  3902 => x"c44b711e",
  3903 => x"fd49d2d9",
  3904 => x"7087f6fb",
  3905 => x"d2d9c44d",
  3906 => x"ecfbfd49",
  3907 => x"c47e7087",
  3908 => x"fd49d2d9",
  3909 => x"7087e2fb",
  3910 => x"05abc44c",
  3911 => x"d9c487c8",
  3912 => x"fbfd49d2",
  3913 => x"487587d3",
  3914 => x"e0c498c7",
  3915 => x"497558f7",
  3916 => x"0299e0c0",
  3917 => x"497487c7",
  3918 => x"71b1c0fc",
  3919 => x"d049754c",
  3920 => x"87c70299",
  3921 => x"c0fc496e",
  3922 => x"c47e71b1",
  3923 => x"48bfebe0",
  3924 => x"e0c4806e",
  3925 => x"497458ef",
  3926 => x"c48909c0",
  3927 => x"48bfefe0",
  3928 => x"e0c48071",
  3929 => x"ef2658f3",
  3930 => x"5e0e87c0",
  3931 => x"0e5d5c5b",
  3932 => x"ff4dd0ff",
  3933 => x"c7c44ad4",
  3934 => x"7dc54bda",
  3935 => x"c37ad5c1",
  3936 => x"c37dc47a",
  3937 => x"7dc57aff",
  3938 => x"c37ad7c1",
  3939 => x"7dc47aff",
  3940 => x"c17dc5c8",
  3941 => x"ffc37ad8",
  3942 => x"ffc34c7a",
  3943 => x"74536a7a",
  3944 => x"718cc149",
  3945 => x"87f20599",
  3946 => x"7dc57dc4",
  3947 => x"c07ad7c1",
  3948 => x"ed7dc47a",
  3949 => x"5e0e87f4",
  3950 => x"0e5d5c5b",
  3951 => x"4dc04b71",
  3952 => x"c04c66d0",
  3953 => x"66d08cf0",
  3954 => x"87edc002",
  3955 => x"028ac34a",
  3956 => x"c087e6c0",
  3957 => x"c1028aed",
  3958 => x"8ac187c4",
  3959 => x"87fec002",
  3960 => x"dbc1028a",
  3961 => x"c1028a87",
  3962 => x"8adf87d6",
  3963 => x"87e1c102",
  3964 => x"c1028ac1",
  3965 => x"d5c287ee",
  3966 => x"029b7387",
  3967 => x"9787cfc2",
  3968 => x"c9c2026b",
  3969 => x"ead9c487",
  3970 => x"b0c248bf",
  3971 => x"58eed9c4",
  3972 => x"7387d9fa",
  3973 => x"f3c8fd49",
  3974 => x"c14d7087",
  3975 => x"1e7487f0",
  3976 => x"f3fe49c0",
  3977 => x"1e7487f4",
  3978 => x"f3fe4973",
  3979 => x"86c887ec",
  3980 => x"c8c14974",
  3981 => x"d3dac491",
  3982 => x"6981c881",
  3983 => x"87cec14d",
  3984 => x"89c24974",
  3985 => x"49731e71",
  3986 => x"87ded7ff",
  3987 => x"fdc086c4",
  3988 => x"cdebc187",
  3989 => x"1e50c348",
  3990 => x"d9fd4973",
  3991 => x"7086c487",
  3992 => x"87eac04d",
  3993 => x"48cdebc1",
  3994 => x"1e7350c3",
  3995 => x"49d0d4c4",
  3996 => x"87ffe7fc",
  3997 => x"987086c4",
  3998 => x"7387d302",
  3999 => x"87eafb49",
  4000 => x"1edac7c4",
  4001 => x"49d0d4c4",
  4002 => x"87ddeefc",
  4003 => x"d9c486c4",
  4004 => x"fd48bfea",
  4005 => x"eed9c498",
  4006 => x"87d0f858",
  4007 => x"c9ea4875",
  4008 => x"1e731e87",
  4009 => x"d9c44bc0",
  4010 => x"78c248ea",
  4011 => x"48c3e0c4",
  4012 => x"d47840c0",
  4013 => x"c878c080",
  4014 => x"c178c380",
  4015 => x"c048cbc1",
  4016 => x"87e8f750",
  4017 => x"48cdebc1",
  4018 => x"c31e50c3",
  4019 => x"fb49e4fc",
  4020 => x"f2c087e4",
  4021 => x"f0fcc31e",
  4022 => x"87dafb49",
  4023 => x"48cdebc1",
  4024 => x"1ec050c1",
  4025 => x"bfccc4c4",
  4026 => x"87cafb49",
  4027 => x"987086cc",
  4028 => x"c387c405",
  4029 => x"c44bfcfc",
  4030 => x"48bfead9",
  4031 => x"d9c498fd",
  4032 => x"e7f658ee",
  4033 => x"87eee887",
  4034 => x"87cef1fd",
  4035 => x"fffd49c1",
  4036 => x"c8c387f5",
  4037 => x"c31ec11e",
  4038 => x"f8e849ff",
  4039 => x"f8487387",
  4040 => x"87cae88e",
  4041 => x"534f4d43",
  4042 => x"20202020",
  4043 => x"004d4152",
  4044 => x"48435241",
  4045 => x"20314549",
  4046 => x"00464448",
  4047 => x"204d4f52",
  4048 => x"64616f6c",
  4049 => x"20676e69",
  4050 => x"6c696166",
  4051 => x"002e6465",
  4052 => x"1e1e731e",
  4053 => x"fefd49c0",
  4054 => x"e7e987ed",
  4055 => x"fe4b7087",
  4056 => x"7387eedf",
  4057 => x"87c8059b",
  4058 => x"87daebfe",
  4059 => x"87e5d3ff",
  4060 => x"ffc1496e",
  4061 => x"486e99ff",
  4062 => x"7e7080c1",
  4063 => x"ff059971",
  4064 => x"e9fd87d2",
  4065 => x"497087cf",
  4066 => x"87d3c6fe",
  4067 => x"2687c5ff",
  4068 => x"7687dbe6",
  4069 => x"0c040605",
  4070 => x"0a830b03",
  4071 => x"07780901",
  4072 => x"0ef77efc",
  4073 => x"25261e16",
  4074 => x"3e3d362e",
  4075 => x"557b4546",
  4076 => x"ecf066ff",
  4077 => x"7cca77fd",
  4078 => x"1d150dff",
  4079 => x"352c2d24",
  4080 => x"4d44433c",
  4081 => x"f15d5b54",
  4082 => x"756cfae9",
  4083 => x"1c14847d",
  4084 => x"342b231b",
  4085 => x"4b423b33",
  4086 => x"6b5a524c",
  4087 => x"12797473",
  4088 => x"21221aff",
  4089 => x"3a31322a",
  4090 => x"594a4941",
  4091 => x"7a7269f5",
  4092 => x"91291158",
  4093 => x"f4f2eb94",
  4094 => x"00da7170",
  4095 => x"f5f2ebf4",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
