
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"e0",x"c4",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"fc",x"e0",x"c4"),
    14 => (x"48",x"f4",x"c6",x"c4"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ea",x"e9"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"1e",x"73",x"1e",x"4f"),
    50 => (x"c0",x"02",x"9a",x"72"),
    51 => (x"48",x"c0",x"87",x"e7"),
    52 => (x"a9",x"72",x"4b",x"c1"),
    53 => (x"72",x"87",x"d1",x"06"),
    54 => (x"87",x"c9",x"06",x"82"),
    55 => (x"a9",x"72",x"83",x"73"),
    56 => (x"c3",x"87",x"f4",x"01"),
    57 => (x"3a",x"b2",x"c1",x"87"),
    58 => (x"89",x"03",x"a9",x"72"),
    59 => (x"c1",x"07",x"80",x"73"),
    60 => (x"f3",x"05",x"2b",x"2a"),
    61 => (x"26",x"4b",x"26",x"87"),
    62 => (x"1e",x"75",x"1e",x"4f"),
    63 => (x"b7",x"71",x"4d",x"c4"),
    64 => (x"b9",x"ff",x"04",x"a1"),
    65 => (x"bd",x"c3",x"81",x"c1"),
    66 => (x"a2",x"b7",x"72",x"07"),
    67 => (x"c1",x"ba",x"ff",x"04"),
    68 => (x"07",x"bd",x"c1",x"82"),
    69 => (x"c1",x"87",x"ee",x"fe"),
    70 => (x"b8",x"ff",x"04",x"2d"),
    71 => (x"2d",x"07",x"80",x"c1"),
    72 => (x"c1",x"b9",x"ff",x"04"),
    73 => (x"4d",x"26",x"07",x"81"),
    74 => (x"71",x"1e",x"4f",x"26"),
    75 => (x"49",x"66",x"c4",x"4a"),
    76 => (x"c8",x"88",x"c1",x"48"),
    77 => (x"99",x"71",x"58",x"a6"),
    78 => (x"12",x"87",x"d4",x"02"),
    79 => (x"08",x"d4",x"ff",x"48"),
    80 => (x"49",x"66",x"c4",x"78"),
    81 => (x"c8",x"88",x"c1",x"48"),
    82 => (x"99",x"71",x"58",x"a6"),
    83 => (x"26",x"87",x"ec",x"05"),
    84 => (x"4a",x"71",x"1e",x"4f"),
    85 => (x"48",x"49",x"66",x"c4"),
    86 => (x"a6",x"c8",x"88",x"c1"),
    87 => (x"02",x"99",x"71",x"58"),
    88 => (x"d4",x"ff",x"87",x"d6"),
    89 => (x"78",x"ff",x"c3",x"48"),
    90 => (x"66",x"c4",x"52",x"68"),
    91 => (x"88",x"c1",x"48",x"49"),
    92 => (x"71",x"58",x"a6",x"c8"),
    93 => (x"87",x"ea",x"05",x"99"),
    94 => (x"73",x"1e",x"4f",x"26"),
    95 => (x"4b",x"d4",x"ff",x"1e"),
    96 => (x"6b",x"7b",x"ff",x"c3"),
    97 => (x"7b",x"ff",x"c3",x"4a"),
    98 => (x"32",x"c8",x"49",x"6b"),
    99 => (x"ff",x"c3",x"b1",x"72"),
   100 => (x"c8",x"4a",x"6b",x"7b"),
   101 => (x"c3",x"b2",x"71",x"31"),
   102 => (x"49",x"6b",x"7b",x"ff"),
   103 => (x"b1",x"72",x"32",x"c8"),
   104 => (x"87",x"c4",x"48",x"71"),
   105 => (x"4c",x"26",x"4d",x"26"),
   106 => (x"4f",x"26",x"4b",x"26"),
   107 => (x"5c",x"5b",x"5e",x"0e"),
   108 => (x"4a",x"71",x"0e",x"5d"),
   109 => (x"72",x"4c",x"d4",x"ff"),
   110 => (x"99",x"ff",x"c3",x"49"),
   111 => (x"c6",x"c4",x"7c",x"71"),
   112 => (x"c8",x"05",x"bf",x"f4"),
   113 => (x"48",x"66",x"d0",x"87"),
   114 => (x"a6",x"d4",x"30",x"c9"),
   115 => (x"49",x"66",x"d0",x"58"),
   116 => (x"ff",x"c3",x"29",x"d8"),
   117 => (x"d0",x"7c",x"71",x"99"),
   118 => (x"29",x"d0",x"49",x"66"),
   119 => (x"71",x"99",x"ff",x"c3"),
   120 => (x"49",x"66",x"d0",x"7c"),
   121 => (x"ff",x"c3",x"29",x"c8"),
   122 => (x"d0",x"7c",x"71",x"99"),
   123 => (x"ff",x"c3",x"49",x"66"),
   124 => (x"72",x"7c",x"71",x"99"),
   125 => (x"c3",x"29",x"d0",x"49"),
   126 => (x"7c",x"71",x"99",x"ff"),
   127 => (x"f0",x"c9",x"4b",x"6c"),
   128 => (x"ff",x"c3",x"4d",x"ff"),
   129 => (x"87",x"d0",x"05",x"ab"),
   130 => (x"6c",x"7c",x"ff",x"c3"),
   131 => (x"02",x"8d",x"c1",x"4b"),
   132 => (x"ff",x"c3",x"87",x"c6"),
   133 => (x"87",x"f0",x"02",x"ab"),
   134 => (x"c7",x"fe",x"48",x"73"),
   135 => (x"49",x"c0",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"81",x"c1",x"78",x"ff"),
   138 => (x"a9",x"b7",x"c8",x"c3"),
   139 => (x"26",x"87",x"f1",x"04"),
   140 => (x"1e",x"73",x"1e",x"4f"),
   141 => (x"f8",x"c4",x"87",x"e7"),
   142 => (x"1e",x"c0",x"4b",x"df"),
   143 => (x"c1",x"f0",x"ff",x"c0"),
   144 => (x"e7",x"fd",x"49",x"f7"),
   145 => (x"c1",x"86",x"c4",x"87"),
   146 => (x"ea",x"c0",x"05",x"a8"),
   147 => (x"48",x"d4",x"ff",x"87"),
   148 => (x"c1",x"78",x"ff",x"c3"),
   149 => (x"c0",x"c0",x"c0",x"c0"),
   150 => (x"e1",x"c0",x"1e",x"c0"),
   151 => (x"49",x"e9",x"c1",x"f0"),
   152 => (x"c4",x"87",x"c9",x"fd"),
   153 => (x"05",x"98",x"70",x"86"),
   154 => (x"d4",x"ff",x"87",x"ca"),
   155 => (x"78",x"ff",x"c3",x"48"),
   156 => (x"87",x"cb",x"48",x"c1"),
   157 => (x"c1",x"87",x"e6",x"fe"),
   158 => (x"fd",x"fe",x"05",x"8b"),
   159 => (x"fc",x"48",x"c0",x"87"),
   160 => (x"73",x"1e",x"87",x"e6"),
   161 => (x"48",x"d4",x"ff",x"1e"),
   162 => (x"d3",x"78",x"ff",x"c3"),
   163 => (x"c0",x"1e",x"c0",x"4b"),
   164 => (x"c1",x"c1",x"f0",x"ff"),
   165 => (x"87",x"d4",x"fc",x"49"),
   166 => (x"98",x"70",x"86",x"c4"),
   167 => (x"ff",x"87",x"ca",x"05"),
   168 => (x"ff",x"c3",x"48",x"d4"),
   169 => (x"cb",x"48",x"c1",x"78"),
   170 => (x"87",x"f1",x"fd",x"87"),
   171 => (x"ff",x"05",x"8b",x"c1"),
   172 => (x"48",x"c0",x"87",x"db"),
   173 => (x"0e",x"87",x"f1",x"fb"),
   174 => (x"0e",x"5c",x"5b",x"5e"),
   175 => (x"fd",x"4c",x"d4",x"ff"),
   176 => (x"ea",x"c6",x"87",x"db"),
   177 => (x"f0",x"e1",x"c0",x"1e"),
   178 => (x"fb",x"49",x"c8",x"c1"),
   179 => (x"86",x"c4",x"87",x"de"),
   180 => (x"c8",x"02",x"a8",x"c1"),
   181 => (x"87",x"ea",x"fe",x"87"),
   182 => (x"e2",x"c1",x"48",x"c0"),
   183 => (x"87",x"da",x"fa",x"87"),
   184 => (x"ff",x"cf",x"49",x"70"),
   185 => (x"ea",x"c6",x"99",x"ff"),
   186 => (x"87",x"c8",x"02",x"a9"),
   187 => (x"c0",x"87",x"d3",x"fe"),
   188 => (x"87",x"cb",x"c1",x"48"),
   189 => (x"c0",x"7c",x"ff",x"c3"),
   190 => (x"f4",x"fc",x"4b",x"f1"),
   191 => (x"02",x"98",x"70",x"87"),
   192 => (x"c0",x"87",x"eb",x"c0"),
   193 => (x"f0",x"ff",x"c0",x"1e"),
   194 => (x"fa",x"49",x"fa",x"c1"),
   195 => (x"86",x"c4",x"87",x"de"),
   196 => (x"d9",x"05",x"98",x"70"),
   197 => (x"7c",x"ff",x"c3",x"87"),
   198 => (x"ff",x"c3",x"49",x"6c"),
   199 => (x"7c",x"7c",x"7c",x"7c"),
   200 => (x"02",x"99",x"c0",x"c1"),
   201 => (x"48",x"c1",x"87",x"c4"),
   202 => (x"48",x"c0",x"87",x"d5"),
   203 => (x"ab",x"c2",x"87",x"d1"),
   204 => (x"c0",x"87",x"c4",x"05"),
   205 => (x"c1",x"87",x"c8",x"48"),
   206 => (x"fd",x"fe",x"05",x"8b"),
   207 => (x"f9",x"48",x"c0",x"87"),
   208 => (x"73",x"1e",x"87",x"e4"),
   209 => (x"f4",x"c6",x"c4",x"1e"),
   210 => (x"c7",x"78",x"c1",x"48"),
   211 => (x"48",x"d0",x"ff",x"4b"),
   212 => (x"c8",x"fb",x"78",x"c2"),
   213 => (x"48",x"d0",x"ff",x"87"),
   214 => (x"1e",x"c0",x"78",x"c3"),
   215 => (x"c1",x"d0",x"e5",x"c0"),
   216 => (x"c7",x"f9",x"49",x"c0"),
   217 => (x"c1",x"86",x"c4",x"87"),
   218 => (x"87",x"c1",x"05",x"a8"),
   219 => (x"05",x"ab",x"c2",x"4b"),
   220 => (x"48",x"c0",x"87",x"c5"),
   221 => (x"c1",x"87",x"f9",x"c0"),
   222 => (x"d0",x"ff",x"05",x"8b"),
   223 => (x"87",x"f7",x"fc",x"87"),
   224 => (x"58",x"f8",x"c6",x"c4"),
   225 => (x"cd",x"05",x"98",x"70"),
   226 => (x"c0",x"1e",x"c1",x"87"),
   227 => (x"d0",x"c1",x"f0",x"ff"),
   228 => (x"87",x"d8",x"f8",x"49"),
   229 => (x"d4",x"ff",x"86",x"c4"),
   230 => (x"78",x"ff",x"c3",x"48"),
   231 => (x"c4",x"87",x"de",x"c4"),
   232 => (x"ff",x"58",x"fc",x"c6"),
   233 => (x"78",x"c2",x"48",x"d0"),
   234 => (x"c3",x"48",x"d4",x"ff"),
   235 => (x"48",x"c1",x"78",x"ff"),
   236 => (x"0e",x"87",x"f5",x"f7"),
   237 => (x"5d",x"5c",x"5b",x"5e"),
   238 => (x"c3",x"4a",x"71",x"0e"),
   239 => (x"d4",x"ff",x"4d",x"ff"),
   240 => (x"ff",x"7c",x"75",x"4c"),
   241 => (x"c3",x"c4",x"48",x"d0"),
   242 => (x"72",x"7c",x"75",x"78"),
   243 => (x"f0",x"ff",x"c0",x"1e"),
   244 => (x"f7",x"49",x"d8",x"c1"),
   245 => (x"86",x"c4",x"87",x"d6"),
   246 => (x"c5",x"02",x"98",x"70"),
   247 => (x"c0",x"48",x"c1",x"87"),
   248 => (x"7c",x"75",x"87",x"f0"),
   249 => (x"c8",x"7c",x"fe",x"c3"),
   250 => (x"66",x"d4",x"1e",x"c0"),
   251 => (x"87",x"fa",x"f4",x"49"),
   252 => (x"7c",x"75",x"86",x"c4"),
   253 => (x"7c",x"75",x"7c",x"75"),
   254 => (x"4b",x"e0",x"da",x"d8"),
   255 => (x"49",x"6c",x"7c",x"75"),
   256 => (x"87",x"c5",x"05",x"99"),
   257 => (x"f3",x"05",x"8b",x"c1"),
   258 => (x"ff",x"7c",x"75",x"87"),
   259 => (x"78",x"c2",x"48",x"d0"),
   260 => (x"cf",x"f6",x"48",x"c0"),
   261 => (x"5b",x"5e",x"0e",x"87"),
   262 => (x"71",x"0e",x"5d",x"5c"),
   263 => (x"c5",x"4c",x"c0",x"4b"),
   264 => (x"4a",x"df",x"cd",x"ee"),
   265 => (x"c3",x"48",x"d4",x"ff"),
   266 => (x"49",x"68",x"78",x"ff"),
   267 => (x"05",x"a9",x"fe",x"c3"),
   268 => (x"70",x"87",x"fd",x"c0"),
   269 => (x"02",x"9b",x"73",x"4d"),
   270 => (x"66",x"d0",x"87",x"cc"),
   271 => (x"f4",x"49",x"73",x"1e"),
   272 => (x"86",x"c4",x"87",x"cf"),
   273 => (x"d0",x"ff",x"87",x"d6"),
   274 => (x"78",x"d1",x"c4",x"48"),
   275 => (x"d0",x"7d",x"ff",x"c3"),
   276 => (x"88",x"c1",x"48",x"66"),
   277 => (x"70",x"58",x"a6",x"d4"),
   278 => (x"87",x"f0",x"05",x"98"),
   279 => (x"c3",x"48",x"d4",x"ff"),
   280 => (x"73",x"78",x"78",x"ff"),
   281 => (x"87",x"c5",x"05",x"9b"),
   282 => (x"d0",x"48",x"d0",x"ff"),
   283 => (x"4c",x"4a",x"c1",x"78"),
   284 => (x"fe",x"05",x"8a",x"c1"),
   285 => (x"48",x"74",x"87",x"ee"),
   286 => (x"1e",x"87",x"e9",x"f4"),
   287 => (x"4a",x"71",x"1e",x"73"),
   288 => (x"d4",x"ff",x"4b",x"c0"),
   289 => (x"78",x"ff",x"c3",x"48"),
   290 => (x"c4",x"48",x"d0",x"ff"),
   291 => (x"d4",x"ff",x"78",x"c3"),
   292 => (x"78",x"ff",x"c3",x"48"),
   293 => (x"ff",x"c0",x"1e",x"72"),
   294 => (x"49",x"d1",x"c1",x"f0"),
   295 => (x"c4",x"87",x"cd",x"f4"),
   296 => (x"05",x"98",x"70",x"86"),
   297 => (x"c0",x"c8",x"87",x"d2"),
   298 => (x"49",x"66",x"cc",x"1e"),
   299 => (x"c4",x"87",x"e6",x"fd"),
   300 => (x"ff",x"4b",x"70",x"86"),
   301 => (x"78",x"c2",x"48",x"d0"),
   302 => (x"eb",x"f3",x"48",x"73"),
   303 => (x"5b",x"5e",x"0e",x"87"),
   304 => (x"c0",x"0e",x"5d",x"5c"),
   305 => (x"f0",x"ff",x"c0",x"1e"),
   306 => (x"f3",x"49",x"c9",x"c1"),
   307 => (x"1e",x"d2",x"87",x"de"),
   308 => (x"49",x"fc",x"c6",x"c4"),
   309 => (x"c8",x"87",x"fe",x"fc"),
   310 => (x"c1",x"4c",x"c0",x"86"),
   311 => (x"ac",x"b7",x"d2",x"84"),
   312 => (x"c4",x"87",x"f8",x"04"),
   313 => (x"bf",x"97",x"fc",x"c6"),
   314 => (x"99",x"c0",x"c3",x"49"),
   315 => (x"05",x"a9",x"c0",x"c1"),
   316 => (x"c4",x"87",x"e7",x"c0"),
   317 => (x"bf",x"97",x"c3",x"c7"),
   318 => (x"c4",x"31",x"d0",x"49"),
   319 => (x"bf",x"97",x"c4",x"c7"),
   320 => (x"72",x"32",x"c8",x"4a"),
   321 => (x"c5",x"c7",x"c4",x"b1"),
   322 => (x"b1",x"4a",x"bf",x"97"),
   323 => (x"ff",x"cf",x"4c",x"71"),
   324 => (x"c1",x"9c",x"ff",x"ff"),
   325 => (x"c1",x"34",x"ca",x"84"),
   326 => (x"c7",x"c4",x"87",x"e7"),
   327 => (x"49",x"bf",x"97",x"c5"),
   328 => (x"99",x"c6",x"31",x"c1"),
   329 => (x"97",x"c6",x"c7",x"c4"),
   330 => (x"b7",x"c7",x"4a",x"bf"),
   331 => (x"c4",x"b1",x"72",x"2a"),
   332 => (x"bf",x"97",x"c1",x"c7"),
   333 => (x"9d",x"cf",x"4d",x"4a"),
   334 => (x"97",x"c2",x"c7",x"c4"),
   335 => (x"9a",x"c3",x"4a",x"bf"),
   336 => (x"c7",x"c4",x"32",x"ca"),
   337 => (x"4b",x"bf",x"97",x"c3"),
   338 => (x"b2",x"73",x"33",x"c2"),
   339 => (x"97",x"c4",x"c7",x"c4"),
   340 => (x"c0",x"c3",x"4b",x"bf"),
   341 => (x"2b",x"b7",x"c6",x"9b"),
   342 => (x"81",x"c2",x"b2",x"73"),
   343 => (x"30",x"71",x"48",x"c1"),
   344 => (x"48",x"c1",x"49",x"70"),
   345 => (x"4d",x"70",x"30",x"75"),
   346 => (x"84",x"c1",x"4c",x"72"),
   347 => (x"c0",x"c8",x"94",x"71"),
   348 => (x"cc",x"06",x"ad",x"b7"),
   349 => (x"b7",x"34",x"c1",x"87"),
   350 => (x"b7",x"c0",x"c8",x"2d"),
   351 => (x"f4",x"ff",x"01",x"ad"),
   352 => (x"f0",x"48",x"74",x"87"),
   353 => (x"5e",x"0e",x"87",x"de"),
   354 => (x"0e",x"5d",x"5c",x"5b"),
   355 => (x"cf",x"c4",x"86",x"f8"),
   356 => (x"78",x"c0",x"48",x"e2"),
   357 => (x"1e",x"da",x"c7",x"c4"),
   358 => (x"de",x"fb",x"49",x"c0"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"ce",x"c9",x"48",x"c0"),
   362 => (x"c1",x"4d",x"c0",x"87"),
   363 => (x"d2",x"fa",x"c0",x"7e"),
   364 => (x"c8",x"c4",x"49",x"bf"),
   365 => (x"c8",x"71",x"4a",x"d0"),
   366 => (x"87",x"ee",x"ea",x"4b"),
   367 => (x"c2",x"05",x"98",x"70"),
   368 => (x"c0",x"7e",x"c0",x"87"),
   369 => (x"49",x"bf",x"ce",x"fa"),
   370 => (x"4a",x"ec",x"c8",x"c4"),
   371 => (x"ea",x"4b",x"c8",x"71"),
   372 => (x"98",x"70",x"87",x"d8"),
   373 => (x"c0",x"87",x"c2",x"05"),
   374 => (x"c0",x"02",x"6e",x"7e"),
   375 => (x"ce",x"c4",x"87",x"fd"),
   376 => (x"c4",x"4d",x"bf",x"e0"),
   377 => (x"bf",x"9f",x"d8",x"cf"),
   378 => (x"d6",x"c5",x"48",x"7e"),
   379 => (x"c7",x"05",x"a8",x"ea"),
   380 => (x"e0",x"ce",x"c4",x"87"),
   381 => (x"87",x"ce",x"4d",x"bf"),
   382 => (x"e9",x"ca",x"48",x"6e"),
   383 => (x"c5",x"02",x"a8",x"d5"),
   384 => (x"c7",x"48",x"c0",x"87"),
   385 => (x"c7",x"c4",x"87",x"f1"),
   386 => (x"49",x"75",x"1e",x"da"),
   387 => (x"c4",x"87",x"ec",x"f9"),
   388 => (x"05",x"98",x"70",x"86"),
   389 => (x"48",x"c0",x"87",x"c5"),
   390 => (x"c0",x"87",x"dc",x"c7"),
   391 => (x"49",x"bf",x"ce",x"fa"),
   392 => (x"4a",x"ec",x"c8",x"c4"),
   393 => (x"e9",x"4b",x"c8",x"71"),
   394 => (x"98",x"70",x"87",x"c0"),
   395 => (x"c4",x"87",x"c8",x"05"),
   396 => (x"c1",x"48",x"e2",x"cf"),
   397 => (x"c0",x"87",x"da",x"78"),
   398 => (x"49",x"bf",x"d2",x"fa"),
   399 => (x"4a",x"d0",x"c8",x"c4"),
   400 => (x"e8",x"4b",x"c8",x"71"),
   401 => (x"98",x"70",x"87",x"e4"),
   402 => (x"87",x"c5",x"c0",x"02"),
   403 => (x"e6",x"c6",x"48",x"c0"),
   404 => (x"d8",x"cf",x"c4",x"87"),
   405 => (x"c1",x"49",x"bf",x"97"),
   406 => (x"c0",x"05",x"a9",x"d5"),
   407 => (x"cf",x"c4",x"87",x"cd"),
   408 => (x"49",x"bf",x"97",x"d9"),
   409 => (x"02",x"a9",x"ea",x"c2"),
   410 => (x"c0",x"87",x"c5",x"c0"),
   411 => (x"87",x"c7",x"c6",x"48"),
   412 => (x"97",x"da",x"c7",x"c4"),
   413 => (x"c3",x"48",x"7e",x"bf"),
   414 => (x"c0",x"02",x"a8",x"e9"),
   415 => (x"48",x"6e",x"87",x"ce"),
   416 => (x"02",x"a8",x"eb",x"c3"),
   417 => (x"c0",x"87",x"c5",x"c0"),
   418 => (x"87",x"eb",x"c5",x"48"),
   419 => (x"97",x"e5",x"c7",x"c4"),
   420 => (x"05",x"99",x"49",x"bf"),
   421 => (x"c4",x"87",x"cc",x"c0"),
   422 => (x"bf",x"97",x"e6",x"c7"),
   423 => (x"02",x"a9",x"c2",x"49"),
   424 => (x"c0",x"87",x"c5",x"c0"),
   425 => (x"87",x"cf",x"c5",x"48"),
   426 => (x"97",x"e7",x"c7",x"c4"),
   427 => (x"cf",x"c4",x"48",x"bf"),
   428 => (x"4c",x"70",x"58",x"de"),
   429 => (x"c4",x"88",x"c1",x"48"),
   430 => (x"c4",x"58",x"e2",x"cf"),
   431 => (x"bf",x"97",x"e8",x"c7"),
   432 => (x"c4",x"81",x"75",x"49"),
   433 => (x"bf",x"97",x"e9",x"c7"),
   434 => (x"72",x"32",x"c8",x"4a"),
   435 => (x"d3",x"c4",x"7e",x"a1"),
   436 => (x"78",x"6e",x"48",x"ef"),
   437 => (x"97",x"ea",x"c7",x"c4"),
   438 => (x"a6",x"c8",x"48",x"bf"),
   439 => (x"e2",x"cf",x"c4",x"58"),
   440 => (x"d4",x"c2",x"02",x"bf"),
   441 => (x"ce",x"fa",x"c0",x"87"),
   442 => (x"c8",x"c4",x"49",x"bf"),
   443 => (x"c8",x"71",x"4a",x"ec"),
   444 => (x"87",x"f6",x"e5",x"4b"),
   445 => (x"c0",x"02",x"98",x"70"),
   446 => (x"48",x"c0",x"87",x"c5"),
   447 => (x"c4",x"87",x"f8",x"c3"),
   448 => (x"4c",x"bf",x"da",x"cf"),
   449 => (x"5c",x"c3",x"d4",x"c4"),
   450 => (x"97",x"ff",x"c7",x"c4"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"fe",x"c7",x"c4"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"97",x"c0",x"c8",x"c4"),
   455 => (x"32",x"d0",x"4a",x"bf"),
   456 => (x"c4",x"49",x"a1",x"72"),
   457 => (x"bf",x"97",x"c1",x"c8"),
   458 => (x"72",x"32",x"d8",x"4a"),
   459 => (x"66",x"c4",x"49",x"a1"),
   460 => (x"ef",x"d3",x"c4",x"91"),
   461 => (x"d3",x"c4",x"81",x"bf"),
   462 => (x"c8",x"c4",x"59",x"f7"),
   463 => (x"4a",x"bf",x"97",x"c7"),
   464 => (x"c8",x"c4",x"32",x"c8"),
   465 => (x"4b",x"bf",x"97",x"c6"),
   466 => (x"c8",x"c4",x"4a",x"a2"),
   467 => (x"4b",x"bf",x"97",x"c8"),
   468 => (x"a2",x"73",x"33",x"d0"),
   469 => (x"c9",x"c8",x"c4",x"4a"),
   470 => (x"cf",x"4b",x"bf",x"97"),
   471 => (x"73",x"33",x"d8",x"9b"),
   472 => (x"d3",x"c4",x"4a",x"a2"),
   473 => (x"d3",x"c4",x"5a",x"fb"),
   474 => (x"c2",x"4a",x"bf",x"f7"),
   475 => (x"c4",x"92",x"74",x"8a"),
   476 => (x"72",x"48",x"fb",x"d3"),
   477 => (x"ca",x"c1",x"78",x"a1"),
   478 => (x"ec",x"c7",x"c4",x"87"),
   479 => (x"c8",x"49",x"bf",x"97"),
   480 => (x"eb",x"c7",x"c4",x"31"),
   481 => (x"a1",x"4a",x"bf",x"97"),
   482 => (x"ea",x"cf",x"c4",x"49"),
   483 => (x"e6",x"cf",x"c4",x"59"),
   484 => (x"31",x"c5",x"49",x"bf"),
   485 => (x"c9",x"81",x"ff",x"c7"),
   486 => (x"c3",x"d4",x"c4",x"29"),
   487 => (x"f1",x"c7",x"c4",x"59"),
   488 => (x"c8",x"4a",x"bf",x"97"),
   489 => (x"f0",x"c7",x"c4",x"32"),
   490 => (x"a2",x"4b",x"bf",x"97"),
   491 => (x"92",x"66",x"c4",x"4a"),
   492 => (x"d3",x"c4",x"82",x"6e"),
   493 => (x"d3",x"c4",x"5a",x"ff"),
   494 => (x"78",x"c0",x"48",x"f7"),
   495 => (x"48",x"f3",x"d3",x"c4"),
   496 => (x"c4",x"78",x"a1",x"72"),
   497 => (x"c4",x"48",x"c3",x"d4"),
   498 => (x"78",x"bf",x"f7",x"d3"),
   499 => (x"48",x"c7",x"d4",x"c4"),
   500 => (x"bf",x"fb",x"d3",x"c4"),
   501 => (x"e2",x"cf",x"c4",x"78"),
   502 => (x"c9",x"c0",x"02",x"bf"),
   503 => (x"c4",x"48",x"74",x"87"),
   504 => (x"c0",x"7e",x"70",x"30"),
   505 => (x"d3",x"c4",x"87",x"c9"),
   506 => (x"c4",x"48",x"bf",x"ff"),
   507 => (x"c4",x"7e",x"70",x"30"),
   508 => (x"6e",x"48",x"e6",x"cf"),
   509 => (x"f8",x"48",x"c1",x"78"),
   510 => (x"26",x"4d",x"26",x"8e"),
   511 => (x"26",x"4b",x"26",x"4c"),
   512 => (x"5b",x"5e",x"0e",x"4f"),
   513 => (x"71",x"0e",x"5d",x"5c"),
   514 => (x"e2",x"cf",x"c4",x"4a"),
   515 => (x"87",x"cb",x"02",x"bf"),
   516 => (x"2b",x"c7",x"4b",x"72"),
   517 => (x"ff",x"c1",x"4c",x"72"),
   518 => (x"72",x"87",x"c9",x"9c"),
   519 => (x"72",x"2b",x"c8",x"4b"),
   520 => (x"9c",x"ff",x"c3",x"4c"),
   521 => (x"bf",x"ef",x"d3",x"c4"),
   522 => (x"ca",x"fa",x"c0",x"83"),
   523 => (x"d9",x"02",x"ab",x"bf"),
   524 => (x"ce",x"fa",x"c0",x"87"),
   525 => (x"da",x"c7",x"c4",x"5b"),
   526 => (x"f0",x"49",x"73",x"1e"),
   527 => (x"86",x"c4",x"87",x"fd"),
   528 => (x"c5",x"05",x"98",x"70"),
   529 => (x"c0",x"48",x"c0",x"87"),
   530 => (x"cf",x"c4",x"87",x"e6"),
   531 => (x"d2",x"02",x"bf",x"e2"),
   532 => (x"c4",x"49",x"74",x"87"),
   533 => (x"da",x"c7",x"c4",x"91"),
   534 => (x"cf",x"4d",x"69",x"81"),
   535 => (x"ff",x"ff",x"ff",x"ff"),
   536 => (x"74",x"87",x"cb",x"9d"),
   537 => (x"c4",x"91",x"c2",x"49"),
   538 => (x"9f",x"81",x"da",x"c7"),
   539 => (x"48",x"75",x"4d",x"69"),
   540 => (x"0e",x"87",x"c6",x"fe"),
   541 => (x"5d",x"5c",x"5b",x"5e"),
   542 => (x"71",x"86",x"f4",x"0e"),
   543 => (x"c5",x"05",x"9c",x"4c"),
   544 => (x"c3",x"48",x"c0",x"87"),
   545 => (x"a4",x"c8",x"87",x"f5"),
   546 => (x"c0",x"48",x"6e",x"7e"),
   547 => (x"02",x"66",x"dc",x"78"),
   548 => (x"66",x"dc",x"87",x"c7"),
   549 => (x"c5",x"05",x"bf",x"97"),
   550 => (x"c3",x"48",x"c0",x"87"),
   551 => (x"1e",x"c0",x"87",x"dd"),
   552 => (x"c9",x"d0",x"49",x"c1"),
   553 => (x"c8",x"86",x"c4",x"87"),
   554 => (x"66",x"c4",x"58",x"a6"),
   555 => (x"87",x"ff",x"c0",x"02"),
   556 => (x"4a",x"ea",x"cf",x"c4"),
   557 => (x"ff",x"49",x"66",x"dc"),
   558 => (x"70",x"87",x"d4",x"de"),
   559 => (x"ee",x"c0",x"02",x"98"),
   560 => (x"4a",x"66",x"c4",x"87"),
   561 => (x"cb",x"49",x"66",x"dc"),
   562 => (x"f7",x"de",x"ff",x"4b"),
   563 => (x"02",x"98",x"70",x"87"),
   564 => (x"1e",x"c0",x"87",x"dd"),
   565 => (x"c4",x"02",x"66",x"c8"),
   566 => (x"c2",x"4d",x"c0",x"87"),
   567 => (x"75",x"4d",x"c1",x"87"),
   568 => (x"87",x"ca",x"cf",x"49"),
   569 => (x"a6",x"c8",x"86",x"c4"),
   570 => (x"05",x"66",x"c4",x"58"),
   571 => (x"c4",x"87",x"c1",x"ff"),
   572 => (x"c4",x"c2",x"02",x"66"),
   573 => (x"81",x"dc",x"49",x"87"),
   574 => (x"78",x"69",x"48",x"6e"),
   575 => (x"da",x"49",x"66",x"c4"),
   576 => (x"4d",x"a4",x"c4",x"81"),
   577 => (x"c4",x"7d",x"69",x"9f"),
   578 => (x"02",x"bf",x"e2",x"cf"),
   579 => (x"66",x"c4",x"87",x"d5"),
   580 => (x"9f",x"81",x"d4",x"49"),
   581 => (x"ff",x"c0",x"49",x"69"),
   582 => (x"48",x"71",x"99",x"ff"),
   583 => (x"a6",x"cc",x"30",x"d0"),
   584 => (x"c8",x"87",x"c5",x"58"),
   585 => (x"78",x"c0",x"48",x"a6"),
   586 => (x"48",x"49",x"66",x"c8"),
   587 => (x"7d",x"70",x"80",x"6d"),
   588 => (x"a4",x"cc",x"7c",x"c0"),
   589 => (x"d0",x"79",x"6d",x"49"),
   590 => (x"79",x"c0",x"49",x"a4"),
   591 => (x"c0",x"48",x"a6",x"c4"),
   592 => (x"4a",x"a4",x"d4",x"78"),
   593 => (x"c8",x"49",x"66",x"c4"),
   594 => (x"49",x"a1",x"72",x"91"),
   595 => (x"79",x"6d",x"41",x"c0"),
   596 => (x"c1",x"48",x"66",x"c4"),
   597 => (x"58",x"a6",x"c8",x"80"),
   598 => (x"04",x"a8",x"b7",x"c6"),
   599 => (x"6e",x"87",x"e2",x"ff"),
   600 => (x"2a",x"c9",x"4a",x"bf"),
   601 => (x"f0",x"c0",x"49",x"72"),
   602 => (x"d8",x"dd",x"ff",x"4a"),
   603 => (x"c1",x"4a",x"70",x"87"),
   604 => (x"72",x"49",x"a4",x"c4"),
   605 => (x"c2",x"48",x"c1",x"79"),
   606 => (x"f4",x"48",x"c0",x"87"),
   607 => (x"87",x"f9",x"f9",x"8e"),
   608 => (x"5c",x"5b",x"5e",x"0e"),
   609 => (x"4c",x"71",x"0e",x"5d"),
   610 => (x"ca",x"c1",x"02",x"9c"),
   611 => (x"49",x"a4",x"c8",x"87"),
   612 => (x"c2",x"c1",x"02",x"69"),
   613 => (x"4a",x"66",x"d0",x"87"),
   614 => (x"d4",x"82",x"49",x"6c"),
   615 => (x"66",x"d0",x"5a",x"a6"),
   616 => (x"cf",x"c4",x"b9",x"4d"),
   617 => (x"ff",x"4a",x"bf",x"de"),
   618 => (x"71",x"99",x"72",x"ba"),
   619 => (x"e4",x"c0",x"02",x"99"),
   620 => (x"4b",x"a4",x"c4",x"87"),
   621 => (x"c8",x"f9",x"49",x"6b"),
   622 => (x"c4",x"7b",x"70",x"87"),
   623 => (x"49",x"bf",x"da",x"cf"),
   624 => (x"7c",x"71",x"81",x"6c"),
   625 => (x"cf",x"c4",x"b9",x"75"),
   626 => (x"ff",x"4a",x"bf",x"de"),
   627 => (x"71",x"99",x"72",x"ba"),
   628 => (x"dc",x"ff",x"05",x"99"),
   629 => (x"f8",x"7c",x"75",x"87"),
   630 => (x"73",x"1e",x"87",x"df"),
   631 => (x"9b",x"4b",x"71",x"1e"),
   632 => (x"c8",x"87",x"c7",x"02"),
   633 => (x"05",x"69",x"49",x"a3"),
   634 => (x"48",x"c0",x"87",x"c5"),
   635 => (x"c4",x"87",x"f7",x"c0"),
   636 => (x"4a",x"bf",x"f3",x"d3"),
   637 => (x"69",x"49",x"a3",x"c4"),
   638 => (x"c4",x"89",x"c2",x"49"),
   639 => (x"91",x"bf",x"da",x"cf"),
   640 => (x"c4",x"4a",x"a2",x"71"),
   641 => (x"49",x"bf",x"de",x"cf"),
   642 => (x"a2",x"71",x"99",x"6b"),
   643 => (x"ce",x"fa",x"c0",x"4a"),
   644 => (x"1e",x"66",x"c8",x"5a"),
   645 => (x"e2",x"e9",x"49",x"72"),
   646 => (x"70",x"86",x"c4",x"87"),
   647 => (x"87",x"c4",x"05",x"98"),
   648 => (x"87",x"c2",x"48",x"c0"),
   649 => (x"d4",x"f7",x"48",x"c1"),
   650 => (x"1e",x"73",x"1e",x"87"),
   651 => (x"02",x"9b",x"4b",x"71"),
   652 => (x"a3",x"c8",x"87",x"c7"),
   653 => (x"c5",x"05",x"69",x"49"),
   654 => (x"c0",x"48",x"c0",x"87"),
   655 => (x"d3",x"c4",x"87",x"f7"),
   656 => (x"c4",x"4a",x"bf",x"f3"),
   657 => (x"49",x"69",x"49",x"a3"),
   658 => (x"cf",x"c4",x"89",x"c2"),
   659 => (x"71",x"91",x"bf",x"da"),
   660 => (x"cf",x"c4",x"4a",x"a2"),
   661 => (x"6b",x"49",x"bf",x"de"),
   662 => (x"4a",x"a2",x"71",x"99"),
   663 => (x"5a",x"ce",x"fa",x"c0"),
   664 => (x"72",x"1e",x"66",x"c8"),
   665 => (x"87",x"cb",x"e5",x"49"),
   666 => (x"98",x"70",x"86",x"c4"),
   667 => (x"c0",x"87",x"c4",x"05"),
   668 => (x"c1",x"87",x"c2",x"48"),
   669 => (x"87",x"c5",x"f6",x"48"),
   670 => (x"5c",x"5b",x"5e",x"0e"),
   671 => (x"86",x"f8",x"0e",x"5d"),
   672 => (x"7e",x"ff",x"4c",x"71"),
   673 => (x"69",x"49",x"a4",x"c8"),
   674 => (x"d4",x"4b",x"c0",x"4d"),
   675 => (x"49",x"73",x"4a",x"a4"),
   676 => (x"a1",x"72",x"91",x"c8"),
   677 => (x"d8",x"49",x"69",x"49"),
   678 => (x"8a",x"71",x"4a",x"66"),
   679 => (x"d8",x"5a",x"a6",x"c8"),
   680 => (x"cc",x"01",x"a9",x"66"),
   681 => (x"b7",x"66",x"c4",x"87"),
   682 => (x"87",x"c5",x"06",x"ad"),
   683 => (x"66",x"c4",x"7e",x"73"),
   684 => (x"c6",x"83",x"c1",x"4d"),
   685 => (x"ff",x"04",x"ab",x"b7"),
   686 => (x"48",x"6e",x"87",x"d1"),
   687 => (x"f8",x"f4",x"8e",x"f8"),
   688 => (x"5b",x"5e",x"0e",x"87"),
   689 => (x"f0",x"0e",x"5d",x"5c"),
   690 => (x"6e",x"7e",x"71",x"86"),
   691 => (x"c4",x"81",x"c8",x"49"),
   692 => (x"78",x"69",x"48",x"a6"),
   693 => (x"78",x"ff",x"80",x"c4"),
   694 => (x"a6",x"d0",x"4d",x"c0"),
   695 => (x"6e",x"4c",x"c0",x"5d"),
   696 => (x"74",x"83",x"d4",x"4b"),
   697 => (x"73",x"92",x"c8",x"4a"),
   698 => (x"66",x"cc",x"4a",x"a2"),
   699 => (x"73",x"91",x"c8",x"49"),
   700 => (x"48",x"6a",x"49",x"a1"),
   701 => (x"49",x"70",x"88",x"69"),
   702 => (x"ad",x"b7",x"c0",x"4d"),
   703 => (x"0d",x"87",x"c2",x"03"),
   704 => (x"ac",x"66",x"cc",x"8d"),
   705 => (x"c4",x"87",x"cd",x"02"),
   706 => (x"03",x"ad",x"b7",x"66"),
   707 => (x"a6",x"cc",x"87",x"c6"),
   708 => (x"5d",x"a6",x"c8",x"5c"),
   709 => (x"b7",x"c6",x"84",x"c1"),
   710 => (x"c2",x"ff",x"04",x"ac"),
   711 => (x"48",x"66",x"cc",x"87"),
   712 => (x"a6",x"d0",x"80",x"c1"),
   713 => (x"a8",x"b7",x"c6",x"58"),
   714 => (x"87",x"f1",x"fe",x"04"),
   715 => (x"f0",x"48",x"66",x"c8"),
   716 => (x"87",x"c5",x"f3",x"8e"),
   717 => (x"5c",x"5b",x"5e",x"0e"),
   718 => (x"86",x"f0",x"0e",x"5d"),
   719 => (x"e0",x"c0",x"4b",x"71"),
   720 => (x"28",x"c9",x"48",x"66"),
   721 => (x"73",x"58",x"a6",x"c8"),
   722 => (x"c6",x"c3",x"02",x"9b"),
   723 => (x"49",x"a3",x"c8",x"87"),
   724 => (x"fe",x"c2",x"02",x"69"),
   725 => (x"de",x"cf",x"c4",x"87"),
   726 => (x"b9",x"ff",x"49",x"bf"),
   727 => (x"66",x"c4",x"48",x"71"),
   728 => (x"58",x"a6",x"cc",x"98"),
   729 => (x"9d",x"6b",x"4d",x"71"),
   730 => (x"6c",x"4c",x"a3",x"c4"),
   731 => (x"ad",x"66",x"c8",x"7e"),
   732 => (x"c4",x"87",x"c6",x"05"),
   733 => (x"c8",x"c2",x"7b",x"66"),
   734 => (x"1e",x"66",x"c8",x"87"),
   735 => (x"f7",x"fb",x"49",x"73"),
   736 => (x"d0",x"86",x"c4",x"87"),
   737 => (x"b7",x"c0",x"58",x"a6"),
   738 => (x"87",x"d1",x"04",x"a8"),
   739 => (x"cc",x"4a",x"a3",x"d4"),
   740 => (x"91",x"c8",x"49",x"66"),
   741 => (x"21",x"49",x"a1",x"72"),
   742 => (x"c7",x"7c",x"69",x"7b"),
   743 => (x"cc",x"7b",x"c0",x"87"),
   744 => (x"7c",x"69",x"49",x"a3"),
   745 => (x"6b",x"48",x"66",x"c4"),
   746 => (x"58",x"a6",x"c8",x"88"),
   747 => (x"49",x"73",x"1e",x"75"),
   748 => (x"c4",x"87",x"c5",x"fb"),
   749 => (x"58",x"a6",x"d0",x"86"),
   750 => (x"49",x"a3",x"c4",x"c1"),
   751 => (x"06",x"ad",x"4a",x"69"),
   752 => (x"cc",x"87",x"f3",x"c0"),
   753 => (x"b7",x"c0",x"48",x"66"),
   754 => (x"e9",x"c0",x"04",x"a8"),
   755 => (x"48",x"a6",x"c8",x"87"),
   756 => (x"cc",x"78",x"a3",x"d4"),
   757 => (x"91",x"c8",x"49",x"66"),
   758 => (x"75",x"81",x"66",x"c8"),
   759 => (x"70",x"88",x"69",x"48"),
   760 => (x"06",x"a9",x"72",x"49"),
   761 => (x"49",x"73",x"87",x"d0"),
   762 => (x"70",x"87",x"d6",x"fb"),
   763 => (x"c8",x"91",x"c8",x"49"),
   764 => (x"41",x"75",x"81",x"66"),
   765 => (x"66",x"c4",x"79",x"6e"),
   766 => (x"49",x"73",x"1e",x"49"),
   767 => (x"c4",x"87",x"c1",x"f6"),
   768 => (x"da",x"c7",x"c4",x"86"),
   769 => (x"f7",x"49",x"73",x"1e"),
   770 => (x"86",x"c4",x"87",x"d0"),
   771 => (x"c0",x"49",x"a3",x"d0"),
   772 => (x"f0",x"79",x"66",x"e0"),
   773 => (x"87",x"e1",x"ef",x"8e"),
   774 => (x"71",x"1e",x"73",x"1e"),
   775 => (x"c0",x"02",x"9b",x"4b"),
   776 => (x"d4",x"c4",x"87",x"e4"),
   777 => (x"4a",x"73",x"5b",x"c7"),
   778 => (x"cf",x"c4",x"8a",x"c2"),
   779 => (x"92",x"49",x"bf",x"da"),
   780 => (x"bf",x"f3",x"d3",x"c4"),
   781 => (x"c4",x"80",x"72",x"48"),
   782 => (x"71",x"58",x"cb",x"d4"),
   783 => (x"c4",x"30",x"c4",x"48"),
   784 => (x"c0",x"58",x"ea",x"cf"),
   785 => (x"d4",x"c4",x"87",x"ed"),
   786 => (x"d3",x"c4",x"48",x"c3"),
   787 => (x"c4",x"78",x"bf",x"f7"),
   788 => (x"c4",x"48",x"c7",x"d4"),
   789 => (x"78",x"bf",x"fb",x"d3"),
   790 => (x"bf",x"e2",x"cf",x"c4"),
   791 => (x"c4",x"87",x"c9",x"02"),
   792 => (x"49",x"bf",x"da",x"cf"),
   793 => (x"87",x"c7",x"31",x"c4"),
   794 => (x"bf",x"ff",x"d3",x"c4"),
   795 => (x"c4",x"31",x"c4",x"49"),
   796 => (x"ee",x"59",x"ea",x"cf"),
   797 => (x"5e",x"0e",x"87",x"c7"),
   798 => (x"71",x"0e",x"5c",x"5b"),
   799 => (x"72",x"4b",x"c0",x"4a"),
   800 => (x"e1",x"c0",x"02",x"9a"),
   801 => (x"49",x"a2",x"da",x"87"),
   802 => (x"c4",x"4b",x"69",x"9f"),
   803 => (x"02",x"bf",x"e2",x"cf"),
   804 => (x"a2",x"d4",x"87",x"cf"),
   805 => (x"49",x"69",x"9f",x"49"),
   806 => (x"ff",x"ff",x"c0",x"4c"),
   807 => (x"c2",x"34",x"d0",x"9c"),
   808 => (x"74",x"4c",x"c0",x"87"),
   809 => (x"49",x"73",x"b3",x"49"),
   810 => (x"ed",x"87",x"ed",x"fd"),
   811 => (x"5e",x"0e",x"87",x"cd"),
   812 => (x"0e",x"5d",x"5c",x"5b"),
   813 => (x"4a",x"71",x"86",x"f4"),
   814 => (x"9a",x"72",x"7e",x"c0"),
   815 => (x"c4",x"87",x"d8",x"02"),
   816 => (x"c0",x"48",x"d6",x"c7"),
   817 => (x"ce",x"c7",x"c4",x"78"),
   818 => (x"c7",x"d4",x"c4",x"48"),
   819 => (x"c7",x"c4",x"78",x"bf"),
   820 => (x"d4",x"c4",x"48",x"d2"),
   821 => (x"c4",x"78",x"bf",x"c3"),
   822 => (x"c0",x"48",x"f7",x"cf"),
   823 => (x"e6",x"cf",x"c4",x"50"),
   824 => (x"c7",x"c4",x"49",x"bf"),
   825 => (x"71",x"4a",x"bf",x"d6"),
   826 => (x"ca",x"c4",x"03",x"aa"),
   827 => (x"cf",x"49",x"72",x"87"),
   828 => (x"ea",x"c0",x"05",x"99"),
   829 => (x"ca",x"fa",x"c0",x"87"),
   830 => (x"ce",x"c7",x"c4",x"48"),
   831 => (x"c7",x"c4",x"78",x"bf"),
   832 => (x"c7",x"c4",x"1e",x"da"),
   833 => (x"c4",x"49",x"bf",x"ce"),
   834 => (x"c1",x"48",x"ce",x"c7"),
   835 => (x"ff",x"71",x"78",x"a1"),
   836 => (x"c4",x"87",x"e8",x"dd"),
   837 => (x"c6",x"fa",x"c0",x"86"),
   838 => (x"da",x"c7",x"c4",x"48"),
   839 => (x"c0",x"87",x"cc",x"78"),
   840 => (x"48",x"bf",x"c6",x"fa"),
   841 => (x"c0",x"80",x"e0",x"c0"),
   842 => (x"c4",x"58",x"ca",x"fa"),
   843 => (x"48",x"bf",x"d6",x"c7"),
   844 => (x"c7",x"c4",x"80",x"c1"),
   845 => (x"86",x"27",x"58",x"da"),
   846 => (x"bf",x"00",x"00",x"0e"),
   847 => (x"9d",x"4d",x"bf",x"97"),
   848 => (x"87",x"e3",x"c2",x"02"),
   849 => (x"02",x"ad",x"e5",x"c3"),
   850 => (x"c0",x"87",x"dc",x"c2"),
   851 => (x"4b",x"bf",x"c6",x"fa"),
   852 => (x"11",x"49",x"a3",x"cb"),
   853 => (x"05",x"ac",x"cf",x"4c"),
   854 => (x"75",x"87",x"d2",x"c1"),
   855 => (x"c1",x"99",x"df",x"49"),
   856 => (x"c4",x"91",x"cd",x"89"),
   857 => (x"c1",x"81",x"ea",x"cf"),
   858 => (x"51",x"12",x"4a",x"a3"),
   859 => (x"12",x"4a",x"a3",x"c3"),
   860 => (x"4a",x"a3",x"c5",x"51"),
   861 => (x"a3",x"c7",x"51",x"12"),
   862 => (x"c9",x"51",x"12",x"4a"),
   863 => (x"51",x"12",x"4a",x"a3"),
   864 => (x"12",x"4a",x"a3",x"ce"),
   865 => (x"4a",x"a3",x"d0",x"51"),
   866 => (x"a3",x"d2",x"51",x"12"),
   867 => (x"d4",x"51",x"12",x"4a"),
   868 => (x"51",x"12",x"4a",x"a3"),
   869 => (x"12",x"4a",x"a3",x"d6"),
   870 => (x"4a",x"a3",x"d8",x"51"),
   871 => (x"a3",x"dc",x"51",x"12"),
   872 => (x"de",x"51",x"12",x"4a"),
   873 => (x"51",x"12",x"4a",x"a3"),
   874 => (x"fa",x"c0",x"7e",x"c1"),
   875 => (x"c8",x"49",x"74",x"87"),
   876 => (x"eb",x"c0",x"05",x"99"),
   877 => (x"d0",x"49",x"74",x"87"),
   878 => (x"87",x"d1",x"05",x"99"),
   879 => (x"c0",x"02",x"66",x"dc"),
   880 => (x"49",x"73",x"87",x"cb"),
   881 => (x"70",x"0f",x"66",x"dc"),
   882 => (x"d3",x"c0",x"02",x"98"),
   883 => (x"c0",x"05",x"6e",x"87"),
   884 => (x"cf",x"c4",x"87",x"c6"),
   885 => (x"50",x"c0",x"48",x"ea"),
   886 => (x"bf",x"c6",x"fa",x"c0"),
   887 => (x"87",x"e1",x"c2",x"48"),
   888 => (x"48",x"f7",x"cf",x"c4"),
   889 => (x"c4",x"7e",x"50",x"c0"),
   890 => (x"49",x"bf",x"e6",x"cf"),
   891 => (x"bf",x"d6",x"c7",x"c4"),
   892 => (x"04",x"aa",x"71",x"4a"),
   893 => (x"c4",x"87",x"f6",x"fb"),
   894 => (x"05",x"bf",x"c7",x"d4"),
   895 => (x"c4",x"87",x"c8",x"c0"),
   896 => (x"02",x"bf",x"e2",x"cf"),
   897 => (x"c4",x"87",x"f8",x"c1"),
   898 => (x"49",x"bf",x"d2",x"c7"),
   899 => (x"70",x"87",x"f2",x"e7"),
   900 => (x"d6",x"c7",x"c4",x"49"),
   901 => (x"48",x"a6",x"c4",x"59"),
   902 => (x"bf",x"d2",x"c7",x"c4"),
   903 => (x"e2",x"cf",x"c4",x"78"),
   904 => (x"d8",x"c0",x"02",x"bf"),
   905 => (x"49",x"66",x"c4",x"87"),
   906 => (x"ff",x"ff",x"ff",x"cf"),
   907 => (x"02",x"a9",x"99",x"f8"),
   908 => (x"c0",x"87",x"c5",x"c0"),
   909 => (x"87",x"e1",x"c0",x"4c"),
   910 => (x"dc",x"c0",x"4c",x"c1"),
   911 => (x"49",x"66",x"c4",x"87"),
   912 => (x"99",x"f8",x"ff",x"cf"),
   913 => (x"c8",x"c0",x"02",x"a9"),
   914 => (x"48",x"a6",x"c8",x"87"),
   915 => (x"c5",x"c0",x"78",x"c0"),
   916 => (x"48",x"a6",x"c8",x"87"),
   917 => (x"66",x"c8",x"78",x"c1"),
   918 => (x"05",x"9c",x"74",x"4c"),
   919 => (x"c4",x"87",x"e0",x"c0"),
   920 => (x"89",x"c2",x"49",x"66"),
   921 => (x"bf",x"da",x"cf",x"c4"),
   922 => (x"d3",x"c4",x"91",x"4a"),
   923 => (x"c4",x"4a",x"bf",x"f3"),
   924 => (x"72",x"48",x"ce",x"c7"),
   925 => (x"c7",x"c4",x"78",x"a1"),
   926 => (x"78",x"c0",x"48",x"d6"),
   927 => (x"c0",x"87",x"de",x"f9"),
   928 => (x"e5",x"8e",x"f4",x"48"),
   929 => (x"00",x"00",x"87",x"f3"),
   930 => (x"ff",x"ff",x"00",x"00"),
   931 => (x"0e",x"96",x"ff",x"ff"),
   932 => (x"0e",x"9f",x"00",x"00"),
   933 => (x"41",x"46",x"00",x"00"),
   934 => (x"20",x"32",x"33",x"54"),
   935 => (x"46",x"00",x"20",x"20"),
   936 => (x"36",x"31",x"54",x"41"),
   937 => (x"00",x"20",x"20",x"20"),
   938 => (x"48",x"d0",x"ff",x"1e"),
   939 => (x"26",x"78",x"e0",x"c0"),
   940 => (x"f8",x"c2",x"1e",x"4f"),
   941 => (x"49",x"70",x"87",x"cd"),
   942 => (x"87",x"c6",x"02",x"99"),
   943 => (x"05",x"a9",x"fb",x"c0"),
   944 => (x"48",x"71",x"87",x"f0"),
   945 => (x"5e",x"0e",x"4f",x"26"),
   946 => (x"71",x"0e",x"5c",x"5b"),
   947 => (x"c2",x"4c",x"c0",x"4b"),
   948 => (x"70",x"87",x"f0",x"f7"),
   949 => (x"c0",x"02",x"99",x"49"),
   950 => (x"ec",x"c0",x"87",x"fa"),
   951 => (x"f3",x"c0",x"02",x"a9"),
   952 => (x"a9",x"fb",x"c0",x"87"),
   953 => (x"87",x"ec",x"c0",x"02"),
   954 => (x"ac",x"b7",x"66",x"cc"),
   955 => (x"d0",x"87",x"c7",x"03"),
   956 => (x"87",x"c2",x"02",x"66"),
   957 => (x"99",x"71",x"53",x"71"),
   958 => (x"c1",x"87",x"c2",x"02"),
   959 => (x"c2",x"f7",x"c2",x"84"),
   960 => (x"99",x"49",x"70",x"87"),
   961 => (x"c0",x"87",x"cd",x"02"),
   962 => (x"c7",x"02",x"a9",x"ec"),
   963 => (x"a9",x"fb",x"c0",x"87"),
   964 => (x"87",x"d4",x"ff",x"05"),
   965 => (x"c3",x"02",x"66",x"d0"),
   966 => (x"7b",x"97",x"c0",x"87"),
   967 => (x"05",x"a9",x"ec",x"c0"),
   968 => (x"4a",x"74",x"87",x"c4"),
   969 => (x"4a",x"74",x"87",x"c5"),
   970 => (x"72",x"8a",x"0a",x"c0"),
   971 => (x"26",x"87",x"c2",x"48"),
   972 => (x"26",x"4c",x"26",x"4d"),
   973 => (x"1e",x"4f",x"26",x"4b"),
   974 => (x"87",x"c7",x"f6",x"c2"),
   975 => (x"c0",x"4a",x"49",x"70"),
   976 => (x"c9",x"04",x"aa",x"f0"),
   977 => (x"aa",x"f9",x"c0",x"87"),
   978 => (x"c0",x"87",x"c3",x"01"),
   979 => (x"c1",x"c1",x"8a",x"f0"),
   980 => (x"87",x"c9",x"04",x"aa"),
   981 => (x"01",x"aa",x"da",x"c1"),
   982 => (x"f7",x"c0",x"87",x"c3"),
   983 => (x"26",x"48",x"72",x"8a"),
   984 => (x"5b",x"5e",x"0e",x"4f"),
   985 => (x"4a",x"71",x"0e",x"5c"),
   986 => (x"72",x"4c",x"d4",x"ff"),
   987 => (x"87",x"e9",x"c0",x"49"),
   988 => (x"02",x"9b",x"4b",x"70"),
   989 => (x"8b",x"c1",x"87",x"c2"),
   990 => (x"c5",x"48",x"d0",x"ff"),
   991 => (x"7c",x"d5",x"c1",x"78"),
   992 => (x"31",x"c6",x"49",x"73"),
   993 => (x"97",x"cd",x"eb",x"c1"),
   994 => (x"71",x"48",x"4a",x"bf"),
   995 => (x"ff",x"7c",x"70",x"b0"),
   996 => (x"78",x"c4",x"48",x"d0"),
   997 => (x"d8",x"fe",x"48",x"73"),
   998 => (x"5b",x"5e",x"0e",x"87"),
   999 => (x"f8",x"0e",x"5d",x"5c"),
  1000 => (x"c0",x"4c",x"71",x"86"),
  1001 => (x"fd",x"f4",x"c2",x"7e"),
  1002 => (x"c1",x"4b",x"c0",x"87"),
  1003 => (x"bf",x"97",x"cb",x"c1"),
  1004 => (x"04",x"a9",x"c0",x"49"),
  1005 => (x"f8",x"fb",x"87",x"cf"),
  1006 => (x"c1",x"83",x"c1",x"87"),
  1007 => (x"bf",x"97",x"cb",x"c1"),
  1008 => (x"f1",x"06",x"ab",x"49"),
  1009 => (x"cb",x"c1",x"c1",x"87"),
  1010 => (x"d0",x"02",x"bf",x"97"),
  1011 => (x"f2",x"f3",x"c2",x"87"),
  1012 => (x"99",x"49",x"70",x"87"),
  1013 => (x"c0",x"87",x"c6",x"02"),
  1014 => (x"f0",x"05",x"a9",x"ec"),
  1015 => (x"c2",x"4b",x"c0",x"87"),
  1016 => (x"70",x"87",x"e0",x"f3"),
  1017 => (x"da",x"f3",x"c2",x"4d"),
  1018 => (x"58",x"a6",x"c8",x"87"),
  1019 => (x"87",x"d3",x"f3",x"c2"),
  1020 => (x"83",x"c1",x"4a",x"70"),
  1021 => (x"97",x"49",x"a4",x"c8"),
  1022 => (x"02",x"ad",x"49",x"69"),
  1023 => (x"ff",x"c0",x"87",x"c7"),
  1024 => (x"e7",x"c0",x"05",x"ad"),
  1025 => (x"49",x"a4",x"c9",x"87"),
  1026 => (x"c4",x"49",x"69",x"97"),
  1027 => (x"c7",x"02",x"a9",x"66"),
  1028 => (x"ff",x"c0",x"48",x"87"),
  1029 => (x"87",x"d4",x"05",x"a8"),
  1030 => (x"97",x"49",x"a4",x"ca"),
  1031 => (x"02",x"aa",x"49",x"69"),
  1032 => (x"ff",x"c0",x"87",x"c6"),
  1033 => (x"87",x"c4",x"05",x"aa"),
  1034 => (x"87",x"d0",x"7e",x"c1"),
  1035 => (x"02",x"ad",x"ec",x"c0"),
  1036 => (x"fb",x"c0",x"87",x"c6"),
  1037 => (x"87",x"c4",x"05",x"ad"),
  1038 => (x"7e",x"c1",x"4b",x"c0"),
  1039 => (x"de",x"fe",x"02",x"6e"),
  1040 => (x"87",x"e4",x"f9",x"87"),
  1041 => (x"8e",x"f8",x"48",x"73"),
  1042 => (x"00",x"87",x"e4",x"fb"),
  1043 => (x"5c",x"5b",x"5e",x"0e"),
  1044 => (x"86",x"f8",x"0e",x"5d"),
  1045 => (x"d4",x"ff",x"4d",x"71"),
  1046 => (x"c4",x"1e",x"75",x"4b"),
  1047 => (x"e0",x"49",x"d0",x"d4"),
  1048 => (x"86",x"c4",x"87",x"d1"),
  1049 => (x"c4",x"02",x"98",x"70"),
  1050 => (x"a6",x"c4",x"87",x"cc"),
  1051 => (x"cf",x"eb",x"c1",x"48"),
  1052 => (x"49",x"75",x"78",x"bf"),
  1053 => (x"ff",x"87",x"ea",x"fb"),
  1054 => (x"78",x"c5",x"48",x"d0"),
  1055 => (x"c0",x"7b",x"d6",x"c1"),
  1056 => (x"49",x"a2",x"75",x"4a"),
  1057 => (x"82",x"c1",x"7b",x"11"),
  1058 => (x"04",x"aa",x"b7",x"cb"),
  1059 => (x"4a",x"cc",x"87",x"f3"),
  1060 => (x"c1",x"7b",x"ff",x"c3"),
  1061 => (x"b7",x"e0",x"c0",x"82"),
  1062 => (x"87",x"f4",x"04",x"aa"),
  1063 => (x"c4",x"48",x"d0",x"ff"),
  1064 => (x"7b",x"ff",x"c3",x"78"),
  1065 => (x"d3",x"c1",x"78",x"c5"),
  1066 => (x"c4",x"7b",x"c1",x"7b"),
  1067 => (x"c0",x"48",x"66",x"78"),
  1068 => (x"c2",x"06",x"a8",x"b7"),
  1069 => (x"d4",x"c4",x"87",x"f0"),
  1070 => (x"c4",x"4c",x"bf",x"d8"),
  1071 => (x"88",x"74",x"48",x"66"),
  1072 => (x"74",x"58",x"a6",x"c8"),
  1073 => (x"f9",x"c1",x"02",x"9c"),
  1074 => (x"da",x"c7",x"c4",x"87"),
  1075 => (x"4d",x"c0",x"c8",x"7e"),
  1076 => (x"ac",x"b7",x"c0",x"8c"),
  1077 => (x"c8",x"87",x"c6",x"03"),
  1078 => (x"c0",x"4d",x"a4",x"c0"),
  1079 => (x"cb",x"d4",x"c4",x"4c"),
  1080 => (x"d0",x"49",x"bf",x"97"),
  1081 => (x"87",x"d1",x"02",x"99"),
  1082 => (x"d4",x"c4",x"1e",x"c0"),
  1083 => (x"e9",x"e3",x"49",x"d0"),
  1084 => (x"70",x"86",x"c4",x"87"),
  1085 => (x"ee",x"c0",x"4a",x"49"),
  1086 => (x"da",x"c7",x"c4",x"87"),
  1087 => (x"d0",x"d4",x"c4",x"1e"),
  1088 => (x"87",x"d6",x"e3",x"49"),
  1089 => (x"49",x"70",x"86",x"c4"),
  1090 => (x"48",x"d0",x"ff",x"4a"),
  1091 => (x"c1",x"78",x"c5",x"c8"),
  1092 => (x"97",x"6e",x"7b",x"d4"),
  1093 => (x"48",x"6e",x"7b",x"bf"),
  1094 => (x"7e",x"70",x"80",x"c1"),
  1095 => (x"ff",x"05",x"8d",x"c1"),
  1096 => (x"d0",x"ff",x"87",x"f0"),
  1097 => (x"72",x"78",x"c4",x"48"),
  1098 => (x"87",x"c5",x"05",x"9a"),
  1099 => (x"c7",x"c1",x"48",x"c0"),
  1100 => (x"c4",x"1e",x"c1",x"87"),
  1101 => (x"e1",x"49",x"d0",x"d4"),
  1102 => (x"86",x"c4",x"87",x"c6"),
  1103 => (x"fe",x"05",x"9c",x"74"),
  1104 => (x"66",x"c4",x"87",x"c7"),
  1105 => (x"a8",x"b7",x"c0",x"48"),
  1106 => (x"c4",x"87",x"d1",x"06"),
  1107 => (x"c0",x"48",x"d0",x"d4"),
  1108 => (x"c0",x"80",x"d0",x"78"),
  1109 => (x"c4",x"80",x"f4",x"78"),
  1110 => (x"78",x"bf",x"dc",x"d4"),
  1111 => (x"c0",x"48",x"66",x"c4"),
  1112 => (x"fd",x"01",x"a8",x"b7"),
  1113 => (x"d0",x"ff",x"87",x"d0"),
  1114 => (x"c1",x"78",x"c5",x"48"),
  1115 => (x"7b",x"c0",x"7b",x"d3"),
  1116 => (x"48",x"c1",x"78",x"c4"),
  1117 => (x"48",x"c0",x"87",x"c2"),
  1118 => (x"4d",x"26",x"8e",x"f8"),
  1119 => (x"4b",x"26",x"4c",x"26"),
  1120 => (x"5e",x"0e",x"4f",x"26"),
  1121 => (x"0e",x"5d",x"5c",x"5b"),
  1122 => (x"c0",x"4b",x"71",x"1e"),
  1123 => (x"04",x"ab",x"4d",x"4c"),
  1124 => (x"c0",x"87",x"e8",x"c0"),
  1125 => (x"75",x"1e",x"d9",x"fe"),
  1126 => (x"87",x"c4",x"02",x"9d"),
  1127 => (x"87",x"c2",x"4a",x"c0"),
  1128 => (x"49",x"72",x"4a",x"c1"),
  1129 => (x"c4",x"87",x"c7",x"ec"),
  1130 => (x"c1",x"7e",x"70",x"86"),
  1131 => (x"c2",x"05",x"6e",x"84"),
  1132 => (x"c1",x"4c",x"73",x"87"),
  1133 => (x"06",x"ac",x"73",x"85"),
  1134 => (x"6e",x"87",x"d8",x"ff"),
  1135 => (x"f9",x"fe",x"26",x"48"),
  1136 => (x"5b",x"5e",x"0e",x"87"),
  1137 => (x"1e",x"0e",x"5d",x"5c"),
  1138 => (x"de",x"49",x"4c",x"71"),
  1139 => (x"ec",x"d5",x"c4",x"91"),
  1140 => (x"97",x"85",x"71",x"4d"),
  1141 => (x"dd",x"c1",x"02",x"6d"),
  1142 => (x"d8",x"d5",x"c4",x"87"),
  1143 => (x"82",x"74",x"4a",x"bf"),
  1144 => (x"dd",x"fe",x"49",x"72"),
  1145 => (x"6e",x"7e",x"70",x"87"),
  1146 => (x"87",x"f3",x"c0",x"02"),
  1147 => (x"4b",x"e0",x"d5",x"c4"),
  1148 => (x"49",x"cb",x"4a",x"6e"),
  1149 => (x"87",x"f0",x"fa",x"fe"),
  1150 => (x"93",x"cb",x"4b",x"74"),
  1151 => (x"83",x"e1",x"eb",x"c1"),
  1152 => (x"c8",x"c1",x"83",x"c4"),
  1153 => (x"49",x"74",x"7b",x"fa"),
  1154 => (x"87",x"cb",x"cf",x"c1"),
  1155 => (x"eb",x"c1",x"7b",x"75"),
  1156 => (x"49",x"bf",x"97",x"ce"),
  1157 => (x"e0",x"d5",x"c4",x"1e"),
  1158 => (x"d9",x"ee",x"c2",x"49"),
  1159 => (x"74",x"86",x"c4",x"87"),
  1160 => (x"f2",x"ce",x"c1",x"49"),
  1161 => (x"c1",x"49",x"c0",x"87"),
  1162 => (x"c4",x"87",x"d1",x"d0"),
  1163 => (x"c0",x"48",x"cc",x"d4"),
  1164 => (x"dd",x"49",x"c1",x"78"),
  1165 => (x"fd",x"26",x"87",x"e1"),
  1166 => (x"6f",x"4c",x"87",x"c0"),
  1167 => (x"6e",x"69",x"64",x"61"),
  1168 => (x"2e",x"2e",x"2e",x"67"),
  1169 => (x"5b",x"5e",x"0e",x"00"),
  1170 => (x"4b",x"71",x"0e",x"5c"),
  1171 => (x"d8",x"d5",x"c4",x"4a"),
  1172 => (x"49",x"72",x"82",x"bf"),
  1173 => (x"70",x"87",x"eb",x"fc"),
  1174 => (x"c4",x"02",x"9c",x"4c"),
  1175 => (x"d5",x"e8",x"49",x"87"),
  1176 => (x"d8",x"d5",x"c4",x"87"),
  1177 => (x"c1",x"78",x"c0",x"48"),
  1178 => (x"87",x"eb",x"dc",x"49"),
  1179 => (x"0e",x"87",x"cd",x"fc"),
  1180 => (x"5d",x"5c",x"5b",x"5e"),
  1181 => (x"c4",x"86",x"f4",x"0e"),
  1182 => (x"c0",x"4d",x"da",x"c7"),
  1183 => (x"48",x"a6",x"c4",x"4c"),
  1184 => (x"d5",x"c4",x"78",x"c0"),
  1185 => (x"c0",x"49",x"bf",x"d8"),
  1186 => (x"c1",x"c1",x"06",x"a9"),
  1187 => (x"da",x"c7",x"c4",x"87"),
  1188 => (x"c0",x"02",x"98",x"48"),
  1189 => (x"fe",x"c0",x"87",x"f8"),
  1190 => (x"66",x"c8",x"1e",x"d9"),
  1191 => (x"c4",x"87",x"c7",x"02"),
  1192 => (x"78",x"c0",x"48",x"a6"),
  1193 => (x"a6",x"c4",x"87",x"c5"),
  1194 => (x"c4",x"78",x"c1",x"48"),
  1195 => (x"fd",x"e7",x"49",x"66"),
  1196 => (x"70",x"86",x"c4",x"87"),
  1197 => (x"c4",x"84",x"c1",x"4d"),
  1198 => (x"80",x"c1",x"48",x"66"),
  1199 => (x"c4",x"58",x"a6",x"c8"),
  1200 => (x"49",x"bf",x"d8",x"d5"),
  1201 => (x"87",x"c6",x"03",x"ac"),
  1202 => (x"ff",x"05",x"9d",x"75"),
  1203 => (x"4c",x"c0",x"87",x"c8"),
  1204 => (x"c3",x"02",x"9d",x"75"),
  1205 => (x"fe",x"c0",x"87",x"e0"),
  1206 => (x"66",x"c8",x"1e",x"d9"),
  1207 => (x"cc",x"87",x"c7",x"02"),
  1208 => (x"78",x"c0",x"48",x"a6"),
  1209 => (x"a6",x"cc",x"87",x"c5"),
  1210 => (x"cc",x"78",x"c1",x"48"),
  1211 => (x"fd",x"e6",x"49",x"66"),
  1212 => (x"70",x"86",x"c4",x"87"),
  1213 => (x"c2",x"02",x"6e",x"7e"),
  1214 => (x"49",x"6e",x"87",x"e9"),
  1215 => (x"69",x"97",x"81",x"cb"),
  1216 => (x"02",x"99",x"d0",x"49"),
  1217 => (x"c1",x"87",x"d6",x"c1"),
  1218 => (x"74",x"4a",x"c5",x"c9"),
  1219 => (x"c1",x"91",x"cb",x"49"),
  1220 => (x"72",x"81",x"e1",x"eb"),
  1221 => (x"c3",x"81",x"c8",x"79"),
  1222 => (x"49",x"74",x"51",x"ff"),
  1223 => (x"d5",x"c4",x"91",x"de"),
  1224 => (x"85",x"71",x"4d",x"ec"),
  1225 => (x"7d",x"97",x"c1",x"c2"),
  1226 => (x"c0",x"49",x"a5",x"c1"),
  1227 => (x"cf",x"c4",x"51",x"e0"),
  1228 => (x"02",x"bf",x"97",x"ea"),
  1229 => (x"84",x"c1",x"87",x"d2"),
  1230 => (x"c4",x"4b",x"a5",x"c2"),
  1231 => (x"db",x"4a",x"ea",x"cf"),
  1232 => (x"e3",x"f5",x"fe",x"49"),
  1233 => (x"87",x"db",x"c1",x"87"),
  1234 => (x"c0",x"49",x"a5",x"cd"),
  1235 => (x"c2",x"84",x"c1",x"51"),
  1236 => (x"4a",x"6e",x"4b",x"a5"),
  1237 => (x"f5",x"fe",x"49",x"cb"),
  1238 => (x"c6",x"c1",x"87",x"ce"),
  1239 => (x"c1",x"c7",x"c1",x"87"),
  1240 => (x"cb",x"49",x"74",x"4a"),
  1241 => (x"e1",x"eb",x"c1",x"91"),
  1242 => (x"c4",x"79",x"72",x"81"),
  1243 => (x"bf",x"97",x"ea",x"cf"),
  1244 => (x"74",x"87",x"d8",x"02"),
  1245 => (x"c1",x"91",x"de",x"49"),
  1246 => (x"ec",x"d5",x"c4",x"84"),
  1247 => (x"c4",x"83",x"71",x"4b"),
  1248 => (x"dd",x"4a",x"ea",x"cf"),
  1249 => (x"df",x"f4",x"fe",x"49"),
  1250 => (x"74",x"87",x"d8",x"87"),
  1251 => (x"c4",x"93",x"de",x"4b"),
  1252 => (x"cb",x"83",x"ec",x"d5"),
  1253 => (x"51",x"c0",x"49",x"a3"),
  1254 => (x"6e",x"73",x"84",x"c1"),
  1255 => (x"fe",x"49",x"cb",x"4a"),
  1256 => (x"c4",x"87",x"c5",x"f4"),
  1257 => (x"80",x"c1",x"48",x"66"),
  1258 => (x"c7",x"58",x"a6",x"c8"),
  1259 => (x"c5",x"c0",x"03",x"ac"),
  1260 => (x"fc",x"05",x"6e",x"87"),
  1261 => (x"48",x"74",x"87",x"e0"),
  1262 => (x"fd",x"f6",x"8e",x"f4"),
  1263 => (x"1e",x"73",x"1e",x"87"),
  1264 => (x"cb",x"49",x"4b",x"71"),
  1265 => (x"e1",x"eb",x"c1",x"91"),
  1266 => (x"4a",x"a1",x"c8",x"81"),
  1267 => (x"48",x"cd",x"eb",x"c1"),
  1268 => (x"a1",x"c9",x"50",x"12"),
  1269 => (x"cb",x"c1",x"c1",x"4a"),
  1270 => (x"ca",x"50",x"12",x"48"),
  1271 => (x"ce",x"eb",x"c1",x"81"),
  1272 => (x"c1",x"50",x"11",x"48"),
  1273 => (x"bf",x"97",x"ce",x"eb"),
  1274 => (x"49",x"c0",x"1e",x"49"),
  1275 => (x"87",x"c6",x"e7",x"c2"),
  1276 => (x"48",x"cc",x"d4",x"c4"),
  1277 => (x"49",x"c1",x"78",x"de"),
  1278 => (x"26",x"87",x"dc",x"d6"),
  1279 => (x"1e",x"87",x"ff",x"f5"),
  1280 => (x"cb",x"49",x"4a",x"71"),
  1281 => (x"e1",x"eb",x"c1",x"91"),
  1282 => (x"11",x"81",x"c8",x"81"),
  1283 => (x"d0",x"d4",x"c4",x"48"),
  1284 => (x"d8",x"d5",x"c4",x"58"),
  1285 => (x"c1",x"78",x"c0",x"48"),
  1286 => (x"87",x"fb",x"d5",x"49"),
  1287 => (x"c0",x"1e",x"4f",x"26"),
  1288 => (x"d7",x"c8",x"c1",x"49"),
  1289 => (x"1e",x"4f",x"26",x"87"),
  1290 => (x"d2",x"02",x"99",x"71"),
  1291 => (x"f6",x"ec",x"c1",x"87"),
  1292 => (x"f7",x"50",x"c0",x"48"),
  1293 => (x"ff",x"cf",x"c1",x"80"),
  1294 => (x"da",x"eb",x"c1",x"40"),
  1295 => (x"c1",x"87",x"ce",x"78"),
  1296 => (x"c1",x"48",x"f2",x"ec"),
  1297 => (x"fc",x"78",x"d3",x"eb"),
  1298 => (x"de",x"d0",x"c1",x"80"),
  1299 => (x"0e",x"4f",x"26",x"78"),
  1300 => (x"0e",x"5c",x"5b",x"5e"),
  1301 => (x"cb",x"4a",x"4c",x"71"),
  1302 => (x"e1",x"eb",x"c1",x"92"),
  1303 => (x"49",x"a2",x"c8",x"82"),
  1304 => (x"97",x"4b",x"a2",x"c9"),
  1305 => (x"97",x"1e",x"4b",x"6b"),
  1306 => (x"ca",x"1e",x"49",x"69"),
  1307 => (x"c0",x"49",x"12",x"82"),
  1308 => (x"c0",x"87",x"d1",x"f3"),
  1309 => (x"87",x"df",x"d4",x"49"),
  1310 => (x"c5",x"c1",x"49",x"74"),
  1311 => (x"8e",x"f8",x"87",x"d9"),
  1312 => (x"1e",x"87",x"f9",x"f3"),
  1313 => (x"4b",x"71",x"1e",x"73"),
  1314 => (x"87",x"c3",x"ff",x"49"),
  1315 => (x"fe",x"fe",x"49",x"73"),
  1316 => (x"87",x"ea",x"f3",x"87"),
  1317 => (x"71",x"1e",x"73",x"1e"),
  1318 => (x"4a",x"a3",x"c6",x"4b"),
  1319 => (x"c1",x"87",x"db",x"02"),
  1320 => (x"87",x"d6",x"02",x"8a"),
  1321 => (x"da",x"c1",x"02",x"8a"),
  1322 => (x"c0",x"02",x"8a",x"87"),
  1323 => (x"02",x"8a",x"87",x"fc"),
  1324 => (x"8a",x"87",x"e1",x"c0"),
  1325 => (x"c1",x"87",x"cb",x"02"),
  1326 => (x"49",x"c7",x"87",x"db"),
  1327 => (x"c1",x"87",x"c0",x"fd"),
  1328 => (x"d5",x"c4",x"87",x"de"),
  1329 => (x"c1",x"02",x"bf",x"d8"),
  1330 => (x"c1",x"48",x"87",x"cb"),
  1331 => (x"dc",x"d5",x"c4",x"88"),
  1332 => (x"87",x"c1",x"c1",x"58"),
  1333 => (x"bf",x"dc",x"d5",x"c4"),
  1334 => (x"87",x"f9",x"c0",x"02"),
  1335 => (x"bf",x"d8",x"d5",x"c4"),
  1336 => (x"c4",x"80",x"c1",x"48"),
  1337 => (x"c0",x"58",x"dc",x"d5"),
  1338 => (x"d5",x"c4",x"87",x"eb"),
  1339 => (x"c6",x"49",x"bf",x"d8"),
  1340 => (x"dc",x"d5",x"c4",x"89"),
  1341 => (x"a9",x"b7",x"c0",x"59"),
  1342 => (x"c4",x"87",x"da",x"03"),
  1343 => (x"c0",x"48",x"d8",x"d5"),
  1344 => (x"c4",x"87",x"d2",x"78"),
  1345 => (x"02",x"bf",x"dc",x"d5"),
  1346 => (x"d5",x"c4",x"87",x"cb"),
  1347 => (x"c6",x"48",x"bf",x"d8"),
  1348 => (x"dc",x"d5",x"c4",x"80"),
  1349 => (x"d1",x"49",x"c0",x"58"),
  1350 => (x"49",x"73",x"87",x"fd"),
  1351 => (x"87",x"f7",x"c2",x"c1"),
  1352 => (x"0e",x"87",x"db",x"f1"),
  1353 => (x"5d",x"5c",x"5b",x"5e"),
  1354 => (x"86",x"d0",x"ff",x"0e"),
  1355 => (x"c8",x"59",x"a6",x"dc"),
  1356 => (x"78",x"c0",x"48",x"a6"),
  1357 => (x"c4",x"c1",x"80",x"c4"),
  1358 => (x"80",x"c4",x"78",x"66"),
  1359 => (x"80",x"c4",x"78",x"c1"),
  1360 => (x"d5",x"c4",x"78",x"c1"),
  1361 => (x"78",x"c1",x"48",x"dc"),
  1362 => (x"bf",x"cc",x"d4",x"c4"),
  1363 => (x"05",x"a8",x"de",x"48"),
  1364 => (x"da",x"f4",x"87",x"cb"),
  1365 => (x"cc",x"49",x"70",x"87"),
  1366 => (x"f9",x"cf",x"59",x"a6"),
  1367 => (x"c5",x"de",x"c2",x"87"),
  1368 => (x"87",x"cd",x"e5",x"87"),
  1369 => (x"87",x"db",x"dd",x"c2"),
  1370 => (x"fb",x"c0",x"4c",x"70"),
  1371 => (x"fb",x"c1",x"02",x"ac"),
  1372 => (x"05",x"66",x"d8",x"87"),
  1373 => (x"c1",x"87",x"ed",x"c1"),
  1374 => (x"c4",x"4a",x"66",x"c0"),
  1375 => (x"72",x"7e",x"6a",x"82"),
  1376 => (x"cb",x"e6",x"c1",x"1e"),
  1377 => (x"49",x"66",x"c4",x"48"),
  1378 => (x"20",x"4a",x"a1",x"c8"),
  1379 => (x"05",x"aa",x"71",x"41"),
  1380 => (x"51",x"10",x"87",x"f9"),
  1381 => (x"c0",x"c1",x"4a",x"26"),
  1382 => (x"ce",x"c1",x"48",x"66"),
  1383 => (x"49",x"6a",x"78",x"fd"),
  1384 => (x"51",x"74",x"81",x"c7"),
  1385 => (x"49",x"66",x"c0",x"c1"),
  1386 => (x"51",x"c1",x"81",x"c8"),
  1387 => (x"49",x"66",x"c0",x"c1"),
  1388 => (x"51",x"c0",x"81",x"c9"),
  1389 => (x"49",x"66",x"c0",x"c1"),
  1390 => (x"51",x"c0",x"81",x"ca"),
  1391 => (x"1e",x"d8",x"1e",x"c1"),
  1392 => (x"81",x"c8",x"49",x"6a"),
  1393 => (x"c8",x"87",x"ff",x"e3"),
  1394 => (x"66",x"c4",x"c1",x"86"),
  1395 => (x"01",x"a8",x"c0",x"48"),
  1396 => (x"a6",x"c8",x"87",x"c7"),
  1397 => (x"ce",x"78",x"c1",x"48"),
  1398 => (x"66",x"c4",x"c1",x"87"),
  1399 => (x"d0",x"88",x"c1",x"48"),
  1400 => (x"87",x"c3",x"58",x"a6"),
  1401 => (x"d0",x"87",x"ca",x"e3"),
  1402 => (x"78",x"c2",x"48",x"a6"),
  1403 => (x"cd",x"02",x"9c",x"74"),
  1404 => (x"66",x"c8",x"87",x"e0"),
  1405 => (x"66",x"c8",x"c1",x"48"),
  1406 => (x"d5",x"cd",x"03",x"a8"),
  1407 => (x"48",x"a6",x"dc",x"87"),
  1408 => (x"80",x"e8",x"78",x"c0"),
  1409 => (x"da",x"c2",x"78",x"c0"),
  1410 => (x"4c",x"70",x"87",x"f9"),
  1411 => (x"05",x"ac",x"d0",x"c1"),
  1412 => (x"c4",x"87",x"da",x"c2"),
  1413 => (x"de",x"e4",x"7e",x"66"),
  1414 => (x"c8",x"49",x"70",x"87"),
  1415 => (x"da",x"c2",x"59",x"a6"),
  1416 => (x"4c",x"70",x"87",x"e1"),
  1417 => (x"05",x"ac",x"ec",x"c0"),
  1418 => (x"c8",x"87",x"ed",x"c1"),
  1419 => (x"91",x"cb",x"49",x"66"),
  1420 => (x"81",x"66",x"c0",x"c1"),
  1421 => (x"6a",x"4a",x"a1",x"c4"),
  1422 => (x"4a",x"a1",x"c8",x"4d"),
  1423 => (x"c1",x"52",x"66",x"c4"),
  1424 => (x"c2",x"79",x"ff",x"cf"),
  1425 => (x"70",x"87",x"fc",x"d9"),
  1426 => (x"d9",x"02",x"9c",x"4c"),
  1427 => (x"ac",x"fb",x"c0",x"87"),
  1428 => (x"74",x"87",x"d3",x"02"),
  1429 => (x"ea",x"d9",x"c2",x"55"),
  1430 => (x"9c",x"4c",x"70",x"87"),
  1431 => (x"c0",x"87",x"c7",x"02"),
  1432 => (x"ff",x"05",x"ac",x"fb"),
  1433 => (x"e0",x"c0",x"87",x"ed"),
  1434 => (x"55",x"c1",x"c2",x"55"),
  1435 => (x"d8",x"7d",x"97",x"c0"),
  1436 => (x"a9",x"6e",x"49",x"66"),
  1437 => (x"c8",x"87",x"db",x"05"),
  1438 => (x"66",x"cc",x"48",x"66"),
  1439 => (x"87",x"ca",x"04",x"a8"),
  1440 => (x"c1",x"48",x"66",x"c8"),
  1441 => (x"58",x"a6",x"cc",x"80"),
  1442 => (x"66",x"cc",x"87",x"c8"),
  1443 => (x"d0",x"88",x"c1",x"48"),
  1444 => (x"d8",x"c2",x"58",x"a6"),
  1445 => (x"4c",x"70",x"87",x"ed"),
  1446 => (x"05",x"ac",x"d0",x"c1"),
  1447 => (x"66",x"d4",x"87",x"c8"),
  1448 => (x"d8",x"80",x"c1",x"48"),
  1449 => (x"d0",x"c1",x"58",x"a6"),
  1450 => (x"e6",x"fd",x"02",x"ac"),
  1451 => (x"a6",x"e0",x"c0",x"87"),
  1452 => (x"78",x"66",x"d8",x"48"),
  1453 => (x"c0",x"48",x"66",x"c4"),
  1454 => (x"05",x"a8",x"66",x"e0"),
  1455 => (x"c0",x"87",x"e5",x"c9"),
  1456 => (x"c0",x"48",x"a6",x"e4"),
  1457 => (x"c0",x"80",x"c4",x"78"),
  1458 => (x"c0",x"48",x"74",x"78"),
  1459 => (x"7e",x"70",x"88",x"fb"),
  1460 => (x"e8",x"c8",x"02",x"6e"),
  1461 => (x"cb",x"48",x"6e",x"87"),
  1462 => (x"6e",x"7e",x"70",x"88"),
  1463 => (x"87",x"ce",x"c1",x"02"),
  1464 => (x"88",x"c9",x"48",x"6e"),
  1465 => (x"02",x"6e",x"7e",x"70"),
  1466 => (x"6e",x"87",x"ea",x"c3"),
  1467 => (x"70",x"88",x"c4",x"48"),
  1468 => (x"ce",x"02",x"6e",x"7e"),
  1469 => (x"c1",x"48",x"6e",x"87"),
  1470 => (x"6e",x"7e",x"70",x"88"),
  1471 => (x"87",x"d5",x"c3",x"02"),
  1472 => (x"dc",x"87",x"f4",x"c7"),
  1473 => (x"f0",x"c0",x"48",x"a6"),
  1474 => (x"f6",x"d6",x"c2",x"78"),
  1475 => (x"c0",x"4c",x"70",x"87"),
  1476 => (x"c0",x"02",x"ac",x"ec"),
  1477 => (x"e0",x"c0",x"87",x"c4"),
  1478 => (x"ec",x"c0",x"5c",x"a6"),
  1479 => (x"cd",x"c0",x"02",x"ac"),
  1480 => (x"de",x"d6",x"c2",x"87"),
  1481 => (x"c0",x"4c",x"70",x"87"),
  1482 => (x"ff",x"05",x"ac",x"ec"),
  1483 => (x"ec",x"c0",x"87",x"f3"),
  1484 => (x"c4",x"c0",x"02",x"ac"),
  1485 => (x"ca",x"d6",x"c2",x"87"),
  1486 => (x"ca",x"1e",x"c0",x"87"),
  1487 => (x"49",x"66",x"d0",x"1e"),
  1488 => (x"c8",x"c1",x"91",x"cb"),
  1489 => (x"80",x"71",x"48",x"66"),
  1490 => (x"c8",x"58",x"a6",x"cc"),
  1491 => (x"80",x"c4",x"48",x"66"),
  1492 => (x"cc",x"58",x"a6",x"d0"),
  1493 => (x"ff",x"49",x"bf",x"66"),
  1494 => (x"c1",x"87",x"eb",x"dd"),
  1495 => (x"d4",x"1e",x"de",x"1e"),
  1496 => (x"ff",x"49",x"bf",x"66"),
  1497 => (x"d0",x"87",x"df",x"dd"),
  1498 => (x"c0",x"49",x"70",x"86"),
  1499 => (x"ec",x"c0",x"89",x"09"),
  1500 => (x"e8",x"c0",x"59",x"a6"),
  1501 => (x"a8",x"c0",x"48",x"66"),
  1502 => (x"87",x"ee",x"c0",x"06"),
  1503 => (x"48",x"66",x"e8",x"c0"),
  1504 => (x"c0",x"03",x"a8",x"dd"),
  1505 => (x"66",x"c4",x"87",x"e4"),
  1506 => (x"e8",x"c0",x"49",x"bf"),
  1507 => (x"e0",x"c0",x"81",x"66"),
  1508 => (x"66",x"e8",x"c0",x"51"),
  1509 => (x"c4",x"81",x"c1",x"49"),
  1510 => (x"c2",x"81",x"bf",x"66"),
  1511 => (x"e8",x"c0",x"51",x"c1"),
  1512 => (x"81",x"c2",x"49",x"66"),
  1513 => (x"81",x"bf",x"66",x"c4"),
  1514 => (x"48",x"6e",x"51",x"c0"),
  1515 => (x"78",x"fd",x"ce",x"c1"),
  1516 => (x"81",x"c8",x"49",x"6e"),
  1517 => (x"6e",x"51",x"66",x"d0"),
  1518 => (x"d4",x"81",x"c9",x"49"),
  1519 => (x"49",x"6e",x"51",x"66"),
  1520 => (x"66",x"dc",x"81",x"ca"),
  1521 => (x"48",x"66",x"d0",x"51"),
  1522 => (x"a6",x"d4",x"80",x"c1"),
  1523 => (x"80",x"d8",x"48",x"58"),
  1524 => (x"e8",x"c4",x"78",x"c1"),
  1525 => (x"de",x"dd",x"ff",x"87"),
  1526 => (x"c0",x"49",x"70",x"87"),
  1527 => (x"ff",x"59",x"a6",x"ec"),
  1528 => (x"70",x"87",x"d4",x"dd"),
  1529 => (x"a6",x"e0",x"c0",x"49"),
  1530 => (x"48",x"66",x"dc",x"59"),
  1531 => (x"05",x"a8",x"ec",x"c0"),
  1532 => (x"dc",x"87",x"ca",x"c0"),
  1533 => (x"e8",x"c0",x"48",x"a6"),
  1534 => (x"c4",x"c0",x"78",x"66"),
  1535 => (x"c2",x"d3",x"c2",x"87"),
  1536 => (x"49",x"66",x"c8",x"87"),
  1537 => (x"c0",x"c1",x"91",x"cb"),
  1538 => (x"80",x"71",x"48",x"66"),
  1539 => (x"4a",x"6e",x"7e",x"70"),
  1540 => (x"49",x"6e",x"82",x"c8"),
  1541 => (x"e8",x"c0",x"81",x"ca"),
  1542 => (x"66",x"dc",x"51",x"66"),
  1543 => (x"c0",x"81",x"c1",x"49"),
  1544 => (x"c1",x"89",x"66",x"e8"),
  1545 => (x"70",x"30",x"71",x"48"),
  1546 => (x"71",x"89",x"c1",x"49"),
  1547 => (x"d9",x"c4",x"7a",x"97"),
  1548 => (x"c0",x"49",x"bf",x"ea"),
  1549 => (x"97",x"29",x"66",x"e8"),
  1550 => (x"71",x"48",x"4a",x"6a"),
  1551 => (x"a6",x"f0",x"c0",x"98"),
  1552 => (x"c4",x"49",x"6e",x"58"),
  1553 => (x"c0",x"4d",x"69",x"81"),
  1554 => (x"c4",x"48",x"66",x"e0"),
  1555 => (x"c0",x"02",x"a8",x"66"),
  1556 => (x"a6",x"c4",x"87",x"c8"),
  1557 => (x"c0",x"78",x"c0",x"48"),
  1558 => (x"a6",x"c4",x"87",x"c5"),
  1559 => (x"c4",x"78",x"c1",x"48"),
  1560 => (x"e0",x"c0",x"1e",x"66"),
  1561 => (x"ff",x"49",x"75",x"1e"),
  1562 => (x"c8",x"87",x"db",x"d9"),
  1563 => (x"c0",x"4c",x"70",x"86"),
  1564 => (x"c1",x"06",x"ac",x"b7"),
  1565 => (x"85",x"74",x"87",x"d4"),
  1566 => (x"74",x"49",x"e0",x"c0"),
  1567 => (x"c1",x"4b",x"75",x"89"),
  1568 => (x"71",x"4a",x"d4",x"e6"),
  1569 => (x"87",x"e0",x"e0",x"fe"),
  1570 => (x"e4",x"c0",x"85",x"c2"),
  1571 => (x"80",x"c1",x"48",x"66"),
  1572 => (x"58",x"a6",x"e8",x"c0"),
  1573 => (x"49",x"66",x"ec",x"c0"),
  1574 => (x"a9",x"70",x"81",x"c1"),
  1575 => (x"87",x"c8",x"c0",x"02"),
  1576 => (x"c0",x"48",x"a6",x"c4"),
  1577 => (x"87",x"c5",x"c0",x"78"),
  1578 => (x"c1",x"48",x"a6",x"c4"),
  1579 => (x"1e",x"66",x"c4",x"78"),
  1580 => (x"c0",x"49",x"a4",x"c2"),
  1581 => (x"88",x"71",x"48",x"e0"),
  1582 => (x"75",x"1e",x"49",x"70"),
  1583 => (x"c5",x"d8",x"ff",x"49"),
  1584 => (x"c0",x"86",x"c8",x"87"),
  1585 => (x"ff",x"01",x"a8",x"b7"),
  1586 => (x"e4",x"c0",x"87",x"c0"),
  1587 => (x"d1",x"c0",x"02",x"66"),
  1588 => (x"c9",x"49",x"6e",x"87"),
  1589 => (x"66",x"e4",x"c0",x"81"),
  1590 => (x"c1",x"48",x"6e",x"51"),
  1591 => (x"c0",x"78",x"cf",x"d1"),
  1592 => (x"49",x"6e",x"87",x"cc"),
  1593 => (x"51",x"c2",x"81",x"c9"),
  1594 => (x"d2",x"c1",x"48",x"6e"),
  1595 => (x"e8",x"c0",x"78",x"c3"),
  1596 => (x"78",x"c1",x"48",x"a6"),
  1597 => (x"ff",x"87",x"c6",x"c0"),
  1598 => (x"70",x"87",x"f6",x"d6"),
  1599 => (x"66",x"e8",x"c0",x"4c"),
  1600 => (x"87",x"f5",x"c0",x"02"),
  1601 => (x"cc",x"48",x"66",x"c8"),
  1602 => (x"c0",x"04",x"a8",x"66"),
  1603 => (x"66",x"c8",x"87",x"cb"),
  1604 => (x"cc",x"80",x"c1",x"48"),
  1605 => (x"e0",x"c0",x"58",x"a6"),
  1606 => (x"48",x"66",x"cc",x"87"),
  1607 => (x"a6",x"d0",x"88",x"c1"),
  1608 => (x"87",x"d5",x"c0",x"58"),
  1609 => (x"05",x"ac",x"c6",x"c1"),
  1610 => (x"d0",x"87",x"c8",x"c0"),
  1611 => (x"80",x"c1",x"48",x"66"),
  1612 => (x"ff",x"58",x"a6",x"d4"),
  1613 => (x"70",x"87",x"fa",x"d5"),
  1614 => (x"48",x"66",x"d4",x"4c"),
  1615 => (x"a6",x"d8",x"80",x"c1"),
  1616 => (x"02",x"9c",x"74",x"58"),
  1617 => (x"c8",x"87",x"cb",x"c0"),
  1618 => (x"c8",x"c1",x"48",x"66"),
  1619 => (x"f2",x"04",x"a8",x"66"),
  1620 => (x"d5",x"ff",x"87",x"eb"),
  1621 => (x"66",x"c8",x"87",x"d2"),
  1622 => (x"03",x"a8",x"c7",x"48"),
  1623 => (x"c4",x"87",x"e5",x"c0"),
  1624 => (x"c0",x"48",x"dc",x"d5"),
  1625 => (x"49",x"66",x"c8",x"78"),
  1626 => (x"c0",x"c1",x"91",x"cb"),
  1627 => (x"a1",x"c4",x"81",x"66"),
  1628 => (x"c0",x"4a",x"6a",x"4a"),
  1629 => (x"66",x"c8",x"79",x"52"),
  1630 => (x"cc",x"80",x"c1",x"48"),
  1631 => (x"a8",x"c7",x"58",x"a6"),
  1632 => (x"87",x"db",x"ff",x"04"),
  1633 => (x"ff",x"8e",x"d0",x"ff"),
  1634 => (x"4c",x"87",x"ef",x"df"),
  1635 => (x"20",x"64",x"61",x"6f"),
  1636 => (x"00",x"20",x"2e",x"2a"),
  1637 => (x"1e",x"00",x"20",x"3a"),
  1638 => (x"4b",x"71",x"1e",x"73"),
  1639 => (x"87",x"c6",x"02",x"9b"),
  1640 => (x"48",x"d8",x"d5",x"c4"),
  1641 => (x"1e",x"c7",x"78",x"c0"),
  1642 => (x"bf",x"d8",x"d5",x"c4"),
  1643 => (x"eb",x"c1",x"1e",x"49"),
  1644 => (x"d4",x"c4",x"1e",x"e1"),
  1645 => (x"ed",x"49",x"bf",x"cc"),
  1646 => (x"86",x"cc",x"87",x"e9"),
  1647 => (x"bf",x"cc",x"d4",x"c4"),
  1648 => (x"87",x"e3",x"e9",x"49"),
  1649 => (x"c8",x"02",x"9b",x"73"),
  1650 => (x"e1",x"eb",x"c1",x"87"),
  1651 => (x"d8",x"f1",x"c0",x"49"),
  1652 => (x"e9",x"de",x"ff",x"87"),
  1653 => (x"1e",x"73",x"1e",x"87"),
  1654 => (x"4b",x"ff",x"c3",x"1e"),
  1655 => (x"fc",x"4a",x"d4",x"ff"),
  1656 => (x"98",x"c1",x"48",x"bf"),
  1657 => (x"02",x"6e",x"7e",x"70"),
  1658 => (x"ff",x"87",x"fb",x"c0"),
  1659 => (x"c1",x"c1",x"48",x"d0"),
  1660 => (x"7a",x"d2",x"c2",x"78"),
  1661 => (x"c7",x"c4",x"7a",x"73"),
  1662 => (x"ff",x"48",x"49",x"db"),
  1663 => (x"73",x"50",x"6a",x"80"),
  1664 => (x"73",x"51",x"6a",x"7a"),
  1665 => (x"6a",x"80",x"c1",x"7a"),
  1666 => (x"6a",x"7a",x"73",x"50"),
  1667 => (x"6a",x"7a",x"73",x"50"),
  1668 => (x"6a",x"7a",x"73",x"49"),
  1669 => (x"6a",x"7a",x"73",x"50"),
  1670 => (x"e4",x"c7",x"c4",x"50"),
  1671 => (x"d0",x"ff",x"59",x"97"),
  1672 => (x"78",x"c0",x"c1",x"48"),
  1673 => (x"c7",x"c4",x"87",x"d7"),
  1674 => (x"ff",x"48",x"49",x"db"),
  1675 => (x"51",x"50",x"c0",x"80"),
  1676 => (x"50",x"c0",x"80",x"c1"),
  1677 => (x"50",x"c1",x"50",x"d9"),
  1678 => (x"c3",x"50",x"e2",x"c0"),
  1679 => (x"e1",x"c7",x"c4",x"50"),
  1680 => (x"f8",x"50",x"c0",x"48"),
  1681 => (x"dc",x"ff",x"26",x"80"),
  1682 => (x"cd",x"1e",x"87",x"f4"),
  1683 => (x"49",x"c1",x"87",x"c1"),
  1684 => (x"fe",x"87",x"c4",x"fd"),
  1685 => (x"70",x"87",x"eb",x"e3"),
  1686 => (x"87",x"cd",x"02",x"98"),
  1687 => (x"87",x"e6",x"ec",x"fe"),
  1688 => (x"c4",x"02",x"98",x"70"),
  1689 => (x"c2",x"4a",x"c1",x"87"),
  1690 => (x"72",x"4a",x"c0",x"87"),
  1691 => (x"87",x"ce",x"05",x"9a"),
  1692 => (x"ea",x"c1",x"1e",x"c0"),
  1693 => (x"fb",x"c0",x"49",x"df"),
  1694 => (x"86",x"c4",x"87",x"d6"),
  1695 => (x"ed",x"c1",x"87",x"fe"),
  1696 => (x"1e",x"c0",x"87",x"e8"),
  1697 => (x"49",x"ea",x"ea",x"c1"),
  1698 => (x"87",x"c4",x"fb",x"c0"),
  1699 => (x"d0",x"c2",x"1e",x"c0"),
  1700 => (x"49",x"70",x"87",x"cf"),
  1701 => (x"87",x"f8",x"fa",x"c0"),
  1702 => (x"f8",x"87",x"ff",x"c2"),
  1703 => (x"53",x"4f",x"26",x"8e"),
  1704 => (x"61",x"66",x"20",x"44"),
  1705 => (x"64",x"65",x"6c",x"69"),
  1706 => (x"6f",x"42",x"00",x"2e"),
  1707 => (x"6e",x"69",x"74",x"6f"),
  1708 => (x"2e",x"2e",x"2e",x"67"),
  1709 => (x"d5",x"c4",x"1e",x"00"),
  1710 => (x"78",x"c0",x"48",x"d8"),
  1711 => (x"48",x"cc",x"d4",x"c4"),
  1712 => (x"c5",x"fe",x"78",x"c0"),
  1713 => (x"c7",x"d2",x"c2",x"87"),
  1714 => (x"26",x"48",x"c0",x"87"),
  1715 => (x"01",x"00",x"00",x"4f"),
  1716 => (x"80",x"00",x"00",x"00"),
  1717 => (x"69",x"78",x"45",x"20"),
  1718 => (x"20",x"80",x"00",x"74"),
  1719 => (x"6b",x"63",x"61",x"42"),
  1720 => (x"00",x"13",x"ff",x"00"),
  1721 => (x"00",x"45",x"6c",x"00"),
  1722 => (x"00",x"00",x"00",x"00"),
  1723 => (x"00",x"00",x"13",x"ff"),
  1724 => (x"00",x"00",x"45",x"8a"),
  1725 => (x"ff",x"00",x"00",x"00"),
  1726 => (x"a8",x"00",x"00",x"13"),
  1727 => (x"00",x"00",x"00",x"45"),
  1728 => (x"13",x"ff",x"00",x"00"),
  1729 => (x"45",x"c6",x"00",x"00"),
  1730 => (x"00",x"00",x"00",x"00"),
  1731 => (x"00",x"13",x"ff",x"00"),
  1732 => (x"00",x"45",x"e4",x"00"),
  1733 => (x"00",x"00",x"00",x"00"),
  1734 => (x"00",x"00",x"13",x"ff"),
  1735 => (x"00",x"00",x"46",x"02"),
  1736 => (x"ff",x"00",x"00",x"00"),
  1737 => (x"20",x"00",x"00",x"13"),
  1738 => (x"00",x"00",x"00",x"46"),
  1739 => (x"13",x"ff",x"00",x"00"),
  1740 => (x"00",x"00",x"00",x"00"),
  1741 => (x"00",x"00",x"00",x"00"),
  1742 => (x"00",x"14",x"94",x"00"),
  1743 => (x"00",x"00",x"00",x"00"),
  1744 => (x"00",x"00",x"00",x"00"),
  1745 => (x"48",x"f0",x"fe",x"1e"),
  1746 => (x"09",x"cd",x"78",x"c0"),
  1747 => (x"4f",x"26",x"09",x"79"),
  1748 => (x"f0",x"fe",x"1e",x"1e"),
  1749 => (x"26",x"48",x"7e",x"bf"),
  1750 => (x"fe",x"1e",x"4f",x"26"),
  1751 => (x"78",x"c1",x"48",x"f0"),
  1752 => (x"fe",x"1e",x"4f",x"26"),
  1753 => (x"78",x"c0",x"48",x"f0"),
  1754 => (x"71",x"1e",x"4f",x"26"),
  1755 => (x"7a",x"97",x"c0",x"4a"),
  1756 => (x"c0",x"49",x"a2",x"c1"),
  1757 => (x"49",x"a2",x"ca",x"51"),
  1758 => (x"a2",x"cb",x"51",x"c0"),
  1759 => (x"26",x"51",x"c0",x"49"),
  1760 => (x"5b",x"5e",x"0e",x"4f"),
  1761 => (x"86",x"f0",x"0e",x"5c"),
  1762 => (x"a4",x"ca",x"4c",x"71"),
  1763 => (x"7e",x"69",x"97",x"49"),
  1764 => (x"97",x"4b",x"a4",x"cb"),
  1765 => (x"a6",x"c8",x"48",x"6b"),
  1766 => (x"cc",x"80",x"c1",x"58"),
  1767 => (x"98",x"c7",x"58",x"a6"),
  1768 => (x"6e",x"58",x"a6",x"d0"),
  1769 => (x"a8",x"66",x"cc",x"48"),
  1770 => (x"97",x"87",x"db",x"05"),
  1771 => (x"6b",x"97",x"7e",x"69"),
  1772 => (x"58",x"a6",x"c8",x"48"),
  1773 => (x"a6",x"cc",x"80",x"c1"),
  1774 => (x"d0",x"98",x"c7",x"58"),
  1775 => (x"48",x"6e",x"58",x"a6"),
  1776 => (x"02",x"a8",x"66",x"cc"),
  1777 => (x"d9",x"fe",x"87",x"e5"),
  1778 => (x"4a",x"a4",x"cc",x"87"),
  1779 => (x"72",x"49",x"6b",x"97"),
  1780 => (x"66",x"dc",x"49",x"a1"),
  1781 => (x"7e",x"6b",x"97",x"51"),
  1782 => (x"80",x"c1",x"48",x"6e"),
  1783 => (x"c7",x"58",x"a6",x"c8"),
  1784 => (x"58",x"a6",x"cc",x"98"),
  1785 => (x"c3",x"7b",x"97",x"70"),
  1786 => (x"ed",x"fd",x"87",x"d2"),
  1787 => (x"c2",x"8e",x"f0",x"87"),
  1788 => (x"26",x"4d",x"26",x"87"),
  1789 => (x"26",x"4b",x"26",x"4c"),
  1790 => (x"5b",x"5e",x"0e",x"4f"),
  1791 => (x"f4",x"0e",x"5d",x"5c"),
  1792 => (x"97",x"4d",x"71",x"86"),
  1793 => (x"a5",x"c1",x"7e",x"6d"),
  1794 => (x"48",x"6c",x"97",x"4c"),
  1795 => (x"6e",x"58",x"a6",x"c8"),
  1796 => (x"a8",x"66",x"c4",x"48"),
  1797 => (x"ff",x"87",x"c5",x"05"),
  1798 => (x"87",x"e6",x"c0",x"48"),
  1799 => (x"c2",x"87",x"c3",x"fd"),
  1800 => (x"6c",x"97",x"49",x"a5"),
  1801 => (x"4b",x"a3",x"71",x"4b"),
  1802 => (x"97",x"4b",x"6b",x"97"),
  1803 => (x"48",x"6e",x"7e",x"6c"),
  1804 => (x"a6",x"c8",x"80",x"c1"),
  1805 => (x"cc",x"98",x"c7",x"58"),
  1806 => (x"97",x"70",x"58",x"a6"),
  1807 => (x"87",x"da",x"fc",x"7c"),
  1808 => (x"8e",x"f4",x"48",x"73"),
  1809 => (x"0e",x"87",x"ea",x"fe"),
  1810 => (x"0e",x"5c",x"5b",x"5e"),
  1811 => (x"4c",x"71",x"86",x"f4"),
  1812 => (x"c3",x"4a",x"66",x"d8"),
  1813 => (x"a4",x"c2",x"9a",x"ff"),
  1814 => (x"49",x"6c",x"97",x"4b"),
  1815 => (x"72",x"49",x"a1",x"73"),
  1816 => (x"7e",x"6c",x"97",x"51"),
  1817 => (x"80",x"c1",x"48",x"6e"),
  1818 => (x"c7",x"58",x"a6",x"c8"),
  1819 => (x"58",x"a6",x"cc",x"98"),
  1820 => (x"8e",x"f4",x"54",x"70"),
  1821 => (x"1e",x"87",x"fc",x"fd"),
  1822 => (x"69",x"97",x"86",x"f0"),
  1823 => (x"4a",x"a1",x"c1",x"7e"),
  1824 => (x"c8",x"48",x"6a",x"97"),
  1825 => (x"48",x"6e",x"58",x"a6"),
  1826 => (x"a8",x"b7",x"66",x"c4"),
  1827 => (x"97",x"87",x"d3",x"04"),
  1828 => (x"6a",x"97",x"7e",x"69"),
  1829 => (x"58",x"a6",x"c8",x"48"),
  1830 => (x"66",x"c4",x"48",x"6e"),
  1831 => (x"58",x"a6",x"cc",x"88"),
  1832 => (x"7e",x"11",x"87",x"d6"),
  1833 => (x"80",x"c8",x"48",x"6e"),
  1834 => (x"48",x"12",x"58",x"a6"),
  1835 => (x"c4",x"58",x"a6",x"cc"),
  1836 => (x"66",x"c8",x"48",x"66"),
  1837 => (x"58",x"a6",x"d0",x"88"),
  1838 => (x"4f",x"26",x"8e",x"f0"),
  1839 => (x"f4",x"1e",x"73",x"1e"),
  1840 => (x"87",x"de",x"fa",x"86"),
  1841 => (x"49",x"4b",x"bf",x"e0"),
  1842 => (x"99",x"c0",x"e0",x"c0"),
  1843 => (x"73",x"87",x"cb",x"02"),
  1844 => (x"fe",x"d8",x"c4",x"1e"),
  1845 => (x"87",x"ef",x"fd",x"49"),
  1846 => (x"49",x"73",x"86",x"c4"),
  1847 => (x"02",x"99",x"c0",x"d0"),
  1848 => (x"c4",x"87",x"c0",x"c1"),
  1849 => (x"bf",x"97",x"c8",x"d9"),
  1850 => (x"c9",x"d9",x"c4",x"7e"),
  1851 => (x"c8",x"48",x"bf",x"97"),
  1852 => (x"48",x"6e",x"58",x"a6"),
  1853 => (x"02",x"a8",x"66",x"c4"),
  1854 => (x"c4",x"87",x"e8",x"c0"),
  1855 => (x"bf",x"97",x"c8",x"d9"),
  1856 => (x"ca",x"d9",x"c4",x"49"),
  1857 => (x"e0",x"48",x"11",x"81"),
  1858 => (x"d9",x"c4",x"78",x"08"),
  1859 => (x"7e",x"bf",x"97",x"c8"),
  1860 => (x"80",x"c1",x"48",x"6e"),
  1861 => (x"c7",x"58",x"a6",x"c8"),
  1862 => (x"58",x"a6",x"cc",x"98"),
  1863 => (x"48",x"c8",x"d9",x"c4"),
  1864 => (x"e4",x"50",x"66",x"c8"),
  1865 => (x"c0",x"49",x"4b",x"bf"),
  1866 => (x"02",x"99",x"c0",x"e0"),
  1867 => (x"1e",x"73",x"87",x"cb"),
  1868 => (x"49",x"d2",x"d9",x"c4"),
  1869 => (x"c4",x"87",x"d0",x"fc"),
  1870 => (x"d0",x"49",x"73",x"86"),
  1871 => (x"c1",x"02",x"99",x"c0"),
  1872 => (x"d9",x"c4",x"87",x"c0"),
  1873 => (x"7e",x"bf",x"97",x"dc"),
  1874 => (x"97",x"dd",x"d9",x"c4"),
  1875 => (x"a6",x"c8",x"48",x"bf"),
  1876 => (x"c4",x"48",x"6e",x"58"),
  1877 => (x"c0",x"02",x"a8",x"66"),
  1878 => (x"d9",x"c4",x"87",x"e8"),
  1879 => (x"49",x"bf",x"97",x"dc"),
  1880 => (x"81",x"de",x"d9",x"c4"),
  1881 => (x"08",x"e4",x"48",x"11"),
  1882 => (x"dc",x"d9",x"c4",x"78"),
  1883 => (x"6e",x"7e",x"bf",x"97"),
  1884 => (x"c8",x"80",x"c1",x"48"),
  1885 => (x"98",x"c7",x"58",x"a6"),
  1886 => (x"c4",x"58",x"a6",x"cc"),
  1887 => (x"c8",x"48",x"dc",x"d9"),
  1888 => (x"cb",x"f7",x"50",x"66"),
  1889 => (x"f7",x"7e",x"70",x"87"),
  1890 => (x"8e",x"f4",x"87",x"d0"),
  1891 => (x"1e",x"87",x"e6",x"f9"),
  1892 => (x"49",x"fe",x"d8",x"c4"),
  1893 => (x"c4",x"87",x"d3",x"f7"),
  1894 => (x"f7",x"49",x"d2",x"d9"),
  1895 => (x"f2",x"c1",x"87",x"cc"),
  1896 => (x"df",x"f6",x"49",x"fc"),
  1897 => (x"87",x"d0",x"c3",x"87"),
  1898 => (x"5e",x"0e",x"4f",x"26"),
  1899 => (x"71",x"0e",x"5c",x"5b"),
  1900 => (x"fe",x"d8",x"c4",x"4c"),
  1901 => (x"87",x"c1",x"f9",x"49"),
  1902 => (x"b7",x"c0",x"4a",x"70"),
  1903 => (x"e3",x"c2",x"04",x"aa"),
  1904 => (x"aa",x"f0",x"c3",x"87"),
  1905 => (x"c1",x"87",x"c9",x"05"),
  1906 => (x"c1",x"48",x"f0",x"f9"),
  1907 => (x"87",x"c4",x"c2",x"78"),
  1908 => (x"05",x"aa",x"e0",x"c3"),
  1909 => (x"f9",x"c1",x"87",x"c9"),
  1910 => (x"78",x"c1",x"48",x"f4"),
  1911 => (x"c1",x"87",x"f5",x"c1"),
  1912 => (x"02",x"bf",x"f4",x"f9"),
  1913 => (x"c0",x"c2",x"87",x"c6"),
  1914 => (x"87",x"c2",x"4b",x"a2"),
  1915 => (x"9c",x"74",x"4b",x"72"),
  1916 => (x"c1",x"87",x"d2",x"05"),
  1917 => (x"1e",x"bf",x"f0",x"f9"),
  1918 => (x"bf",x"f4",x"f9",x"c1"),
  1919 => (x"c1",x"49",x"72",x"1e"),
  1920 => (x"c8",x"87",x"d1",x"f8"),
  1921 => (x"f0",x"f9",x"c1",x"86"),
  1922 => (x"e0",x"c0",x"02",x"bf"),
  1923 => (x"c4",x"49",x"73",x"87"),
  1924 => (x"c1",x"91",x"29",x"b7"),
  1925 => (x"73",x"81",x"c7",x"fb"),
  1926 => (x"c2",x"9a",x"cf",x"4a"),
  1927 => (x"72",x"48",x"c1",x"92"),
  1928 => (x"ff",x"4a",x"70",x"30"),
  1929 => (x"69",x"48",x"72",x"ba"),
  1930 => (x"db",x"79",x"70",x"98"),
  1931 => (x"c4",x"49",x"73",x"87"),
  1932 => (x"c1",x"91",x"29",x"b7"),
  1933 => (x"73",x"81",x"c7",x"fb"),
  1934 => (x"c2",x"9a",x"cf",x"4a"),
  1935 => (x"72",x"48",x"c3",x"92"),
  1936 => (x"48",x"4a",x"70",x"30"),
  1937 => (x"79",x"70",x"b0",x"69"),
  1938 => (x"48",x"f4",x"f9",x"c1"),
  1939 => (x"f9",x"c1",x"78",x"c0"),
  1940 => (x"78",x"c0",x"48",x"f0"),
  1941 => (x"49",x"fe",x"d8",x"c4"),
  1942 => (x"70",x"87",x"de",x"f6"),
  1943 => (x"aa",x"b7",x"c0",x"4a"),
  1944 => (x"87",x"dd",x"fd",x"03"),
  1945 => (x"87",x"c2",x"48",x"c0"),
  1946 => (x"4c",x"26",x"4d",x"26"),
  1947 => (x"4f",x"26",x"4b",x"26"),
  1948 => (x"00",x"00",x"00",x"00"),
  1949 => (x"00",x"00",x"00",x"00"),
  1950 => (x"72",x"4a",x"c0",x"1e"),
  1951 => (x"c1",x"91",x"c4",x"49"),
  1952 => (x"c0",x"81",x"c7",x"fb"),
  1953 => (x"d0",x"82",x"c1",x"79"),
  1954 => (x"ee",x"04",x"aa",x"b7"),
  1955 => (x"0e",x"4f",x"26",x"87"),
  1956 => (x"5d",x"5c",x"5b",x"5e"),
  1957 => (x"f3",x"4d",x"71",x"0e"),
  1958 => (x"4a",x"75",x"87",x"c8"),
  1959 => (x"92",x"2a",x"b7",x"c4"),
  1960 => (x"82",x"c7",x"fb",x"c1"),
  1961 => (x"9c",x"cf",x"4c",x"75"),
  1962 => (x"49",x"6a",x"94",x"c2"),
  1963 => (x"c3",x"2b",x"74",x"4b"),
  1964 => (x"74",x"48",x"c2",x"9b"),
  1965 => (x"ff",x"4c",x"70",x"30"),
  1966 => (x"71",x"48",x"74",x"bc"),
  1967 => (x"f2",x"7a",x"70",x"98"),
  1968 => (x"48",x"73",x"87",x"d8"),
  1969 => (x"00",x"87",x"e1",x"fe"),
  1970 => (x"00",x"00",x"00",x"00"),
  1971 => (x"00",x"00",x"00",x"00"),
  1972 => (x"00",x"00",x"00",x"00"),
  1973 => (x"00",x"00",x"00",x"00"),
  1974 => (x"00",x"00",x"00",x"00"),
  1975 => (x"00",x"00",x"00",x"00"),
  1976 => (x"00",x"00",x"00",x"00"),
  1977 => (x"00",x"00",x"00",x"00"),
  1978 => (x"00",x"00",x"00",x"00"),
  1979 => (x"00",x"00",x"00",x"00"),
  1980 => (x"00",x"00",x"00",x"00"),
  1981 => (x"00",x"00",x"00",x"00"),
  1982 => (x"00",x"00",x"00",x"00"),
  1983 => (x"00",x"00",x"00",x"00"),
  1984 => (x"00",x"00",x"00",x"00"),
  1985 => (x"0e",x"00",x"00",x"00"),
  1986 => (x"5d",x"5c",x"5b",x"5e"),
  1987 => (x"9a",x"4a",x"71",x"0e"),
  1988 => (x"c2",x"87",x"c6",x"02"),
  1989 => (x"c0",x"48",x"e8",x"c2"),
  1990 => (x"e8",x"c2",x"c2",x"78"),
  1991 => (x"c6",x"c1",x"05",x"bf"),
  1992 => (x"d2",x"d9",x"c4",x"87"),
  1993 => (x"87",x"d1",x"f3",x"49"),
  1994 => (x"04",x"a8",x"b7",x"c0"),
  1995 => (x"d9",x"c4",x"87",x"cd"),
  1996 => (x"c4",x"f3",x"49",x"d2"),
  1997 => (x"a8",x"b7",x"c0",x"87"),
  1998 => (x"c2",x"87",x"f3",x"03"),
  1999 => (x"49",x"bf",x"e8",x"c2"),
  2000 => (x"48",x"e8",x"c2",x"c2"),
  2001 => (x"c2",x"78",x"a1",x"c1"),
  2002 => (x"11",x"81",x"f8",x"c2"),
  2003 => (x"f0",x"c2",x"c2",x"48"),
  2004 => (x"f0",x"c2",x"c2",x"58"),
  2005 => (x"c0",x"78",x"c0",x"48"),
  2006 => (x"e9",x"c0",x"49",x"f2"),
  2007 => (x"49",x"70",x"87",x"cf"),
  2008 => (x"59",x"ea",x"d9",x"c4"),
  2009 => (x"c2",x"87",x"f9",x"c4"),
  2010 => (x"02",x"bf",x"f0",x"c2"),
  2011 => (x"c4",x"87",x"f2",x"c1"),
  2012 => (x"f2",x"49",x"d2",x"d9"),
  2013 => (x"b7",x"c0",x"87",x"c3"),
  2014 => (x"87",x"cd",x"04",x"a8"),
  2015 => (x"bf",x"f0",x"c2",x"c2"),
  2016 => (x"c2",x"88",x"c1",x"48"),
  2017 => (x"db",x"58",x"f4",x"c2"),
  2018 => (x"e6",x"d9",x"c4",x"87"),
  2019 => (x"e8",x"c0",x"49",x"bf"),
  2020 => (x"98",x"70",x"87",x"e7"),
  2021 => (x"c4",x"87",x"cd",x"02"),
  2022 => (x"ef",x"49",x"d2",x"d9"),
  2023 => (x"c2",x"c2",x"87",x"cc"),
  2024 => (x"78",x"c0",x"48",x"e8"),
  2025 => (x"bf",x"ec",x"c2",x"c2"),
  2026 => (x"87",x"f4",x"c3",x"05"),
  2027 => (x"bf",x"f0",x"c2",x"c2"),
  2028 => (x"87",x"ec",x"c3",x"05"),
  2029 => (x"bf",x"e8",x"c2",x"c2"),
  2030 => (x"e8",x"c2",x"c2",x"49"),
  2031 => (x"78",x"a1",x"c1",x"48"),
  2032 => (x"81",x"f8",x"c2",x"c2"),
  2033 => (x"c2",x"49",x"4b",x"11"),
  2034 => (x"c0",x"02",x"99",x"c0"),
  2035 => (x"48",x"73",x"87",x"cc"),
  2036 => (x"c2",x"98",x"ff",x"c1"),
  2037 => (x"c3",x"58",x"f4",x"c2"),
  2038 => (x"c2",x"c2",x"87",x"c6"),
  2039 => (x"ff",x"c2",x"5b",x"f0"),
  2040 => (x"ec",x"c2",x"c2",x"87"),
  2041 => (x"db",x"c1",x"02",x"bf"),
  2042 => (x"e6",x"d9",x"c4",x"87"),
  2043 => (x"e7",x"c0",x"49",x"bf"),
  2044 => (x"98",x"70",x"87",x"c7"),
  2045 => (x"87",x"e8",x"c2",x"02"),
  2046 => (x"bf",x"e8",x"c2",x"c2"),
  2047 => (x"e8",x"c2",x"c2",x"49"),
  2048 => (x"78",x"a1",x"c1",x"48"),
  2049 => (x"81",x"f8",x"c2",x"c2"),
  2050 => (x"1e",x"49",x"69",x"97"),
  2051 => (x"49",x"d2",x"d9",x"c4"),
  2052 => (x"c4",x"87",x"ee",x"ed"),
  2053 => (x"ec",x"c2",x"c2",x"86"),
  2054 => (x"89",x"c1",x"49",x"bf"),
  2055 => (x"59",x"f0",x"c2",x"c2"),
  2056 => (x"48",x"f0",x"c2",x"c2"),
  2057 => (x"99",x"71",x"78",x"c1"),
  2058 => (x"87",x"c6",x"c0",x"02"),
  2059 => (x"c0",x"4c",x"f2",x"c0"),
  2060 => (x"dc",x"d7",x"87",x"c3"),
  2061 => (x"c0",x"49",x"74",x"4c"),
  2062 => (x"70",x"87",x"f2",x"e5"),
  2063 => (x"ea",x"d9",x"c4",x"49"),
  2064 => (x"87",x"dc",x"c1",x"59"),
  2065 => (x"49",x"d2",x"d9",x"c4"),
  2066 => (x"70",x"87",x"ec",x"f0"),
  2067 => (x"c0",x"02",x"9b",x"4b"),
  2068 => (x"c2",x"c2",x"87",x"ee"),
  2069 => (x"ab",x"b7",x"bf",x"f4"),
  2070 => (x"87",x"e4",x"c0",x"03"),
  2071 => (x"bf",x"e6",x"d9",x"c4"),
  2072 => (x"d4",x"e5",x"c0",x"49"),
  2073 => (x"02",x"98",x"70",x"87"),
  2074 => (x"c7",x"87",x"f5",x"c0"),
  2075 => (x"f4",x"c2",x"c2",x"48"),
  2076 => (x"c2",x"c2",x"88",x"bf"),
  2077 => (x"d9",x"c4",x"58",x"f8"),
  2078 => (x"ed",x"eb",x"49",x"d2"),
  2079 => (x"87",x"e0",x"c0",x"87"),
  2080 => (x"c0",x"49",x"dc",x"d7"),
  2081 => (x"70",x"87",x"e6",x"e4"),
  2082 => (x"ea",x"d9",x"c4",x"49"),
  2083 => (x"f4",x"c2",x"c2",x"59"),
  2084 => (x"ab",x"b7",x"4a",x"bf"),
  2085 => (x"87",x"c8",x"c0",x"04"),
  2086 => (x"d5",x"f1",x"c1",x"49"),
  2087 => (x"87",x"e4",x"fe",x"87"),
  2088 => (x"4c",x"26",x"4d",x"26"),
  2089 => (x"4f",x"26",x"4b",x"26"),
  2090 => (x"00",x"00",x"00",x"00"),
  2091 => (x"00",x"00",x"00",x"00"),
  2092 => (x"00",x"00",x"00",x"00"),
  2093 => (x"00",x"00",x"00",x"04"),
  2094 => (x"08",x"82",x"ff",x"01"),
  2095 => (x"64",x"f3",x"c8",x"f3"),
  2096 => (x"01",x"f2",x"50",x"f3"),
  2097 => (x"00",x"f4",x"01",x"81"),
  2098 => (x"48",x"d0",x"ff",x"1e"),
  2099 => (x"71",x"78",x"e1",x"c8"),
  2100 => (x"08",x"d4",x"ff",x"48"),
  2101 => (x"1e",x"4f",x"26",x"78"),
  2102 => (x"c8",x"48",x"d0",x"ff"),
  2103 => (x"48",x"71",x"78",x"e1"),
  2104 => (x"78",x"08",x"d4",x"ff"),
  2105 => (x"ff",x"48",x"66",x"c4"),
  2106 => (x"26",x"78",x"08",x"d4"),
  2107 => (x"4a",x"71",x"1e",x"4f"),
  2108 => (x"1e",x"49",x"66",x"c4"),
  2109 => (x"de",x"ff",x"49",x"72"),
  2110 => (x"48",x"d0",x"ff",x"87"),
  2111 => (x"26",x"78",x"e0",x"c0"),
  2112 => (x"73",x"1e",x"4f",x"26"),
  2113 => (x"c8",x"4b",x"71",x"1e"),
  2114 => (x"73",x"1e",x"49",x"66"),
  2115 => (x"a2",x"e0",x"c1",x"4a"),
  2116 => (x"87",x"d9",x"ff",x"49"),
  2117 => (x"26",x"87",x"c4",x"26"),
  2118 => (x"26",x"4c",x"26",x"4d"),
  2119 => (x"1e",x"4f",x"26",x"4b"),
  2120 => (x"4b",x"71",x"1e",x"73"),
  2121 => (x"fe",x"49",x"e2",x"c0"),
  2122 => (x"4a",x"c7",x"87",x"de"),
  2123 => (x"d4",x"ff",x"48",x"13"),
  2124 => (x"49",x"72",x"78",x"08"),
  2125 => (x"99",x"71",x"8a",x"c1"),
  2126 => (x"ff",x"87",x"f1",x"05"),
  2127 => (x"e0",x"c0",x"48",x"d0"),
  2128 => (x"87",x"d7",x"ff",x"78"),
  2129 => (x"5c",x"5b",x"5e",x"0e"),
  2130 => (x"4c",x"71",x"0e",x"5d"),
  2131 => (x"bf",x"ea",x"d9",x"c4"),
  2132 => (x"2b",x"74",x"4b",x"4d"),
  2133 => (x"c1",x"9b",x"66",x"d0"),
  2134 => (x"ab",x"66",x"d4",x"83"),
  2135 => (x"c0",x"87",x"c2",x"04"),
  2136 => (x"d0",x"4a",x"74",x"4b"),
  2137 => (x"31",x"72",x"49",x"66"),
  2138 => (x"99",x"75",x"b9",x"ff"),
  2139 => (x"30",x"72",x"48",x"73"),
  2140 => (x"71",x"48",x"4a",x"70"),
  2141 => (x"ee",x"d9",x"c4",x"b0"),
  2142 => (x"ef",x"ec",x"c1",x"58"),
  2143 => (x"26",x"4d",x"26",x"87"),
  2144 => (x"26",x"4b",x"26",x"4c"),
  2145 => (x"d0",x"ff",x"1e",x"4f"),
  2146 => (x"78",x"c9",x"c8",x"48"),
  2147 => (x"d4",x"ff",x"48",x"71"),
  2148 => (x"4f",x"26",x"78",x"08"),
  2149 => (x"49",x"4a",x"71",x"1e"),
  2150 => (x"d0",x"ff",x"87",x"eb"),
  2151 => (x"26",x"78",x"c8",x"48"),
  2152 => (x"1e",x"73",x"1e",x"4f"),
  2153 => (x"d9",x"c4",x"4b",x"71"),
  2154 => (x"c3",x"02",x"bf",x"fa"),
  2155 => (x"87",x"eb",x"c2",x"87"),
  2156 => (x"c8",x"48",x"d0",x"ff"),
  2157 => (x"49",x"73",x"78",x"c9"),
  2158 => (x"ff",x"b1",x"e0",x"c0"),
  2159 => (x"78",x"71",x"48",x"d4"),
  2160 => (x"48",x"ee",x"d9",x"c4"),
  2161 => (x"66",x"c8",x"78",x"c0"),
  2162 => (x"c3",x"87",x"c5",x"02"),
  2163 => (x"87",x"c2",x"49",x"ff"),
  2164 => (x"d9",x"c4",x"49",x"c0"),
  2165 => (x"66",x"cc",x"59",x"f6"),
  2166 => (x"c5",x"87",x"c6",x"02"),
  2167 => (x"c4",x"4a",x"d5",x"d5"),
  2168 => (x"ff",x"ff",x"cf",x"87"),
  2169 => (x"fa",x"d9",x"c4",x"4a"),
  2170 => (x"fa",x"d9",x"c4",x"5a"),
  2171 => (x"c4",x"78",x"c1",x"48"),
  2172 => (x"26",x"4d",x"26",x"87"),
  2173 => (x"26",x"4b",x"26",x"4c"),
  2174 => (x"5b",x"5e",x"0e",x"4f"),
  2175 => (x"71",x"0e",x"5d",x"5c"),
  2176 => (x"f6",x"d9",x"c4",x"4a"),
  2177 => (x"9a",x"72",x"4c",x"bf"),
  2178 => (x"49",x"87",x"cb",x"02"),
  2179 => (x"c6",x"c2",x"91",x"c8"),
  2180 => (x"83",x"71",x"4b",x"d7"),
  2181 => (x"ca",x"c2",x"87",x"c4"),
  2182 => (x"4d",x"c0",x"4b",x"d7"),
  2183 => (x"99",x"74",x"49",x"13"),
  2184 => (x"bf",x"f2",x"d9",x"c4"),
  2185 => (x"48",x"d4",x"ff",x"b9"),
  2186 => (x"b7",x"c1",x"78",x"71"),
  2187 => (x"b7",x"c8",x"85",x"2c"),
  2188 => (x"87",x"e8",x"04",x"ad"),
  2189 => (x"bf",x"ee",x"d9",x"c4"),
  2190 => (x"c4",x"80",x"c8",x"48"),
  2191 => (x"fe",x"58",x"f2",x"d9"),
  2192 => (x"73",x"1e",x"87",x"ef"),
  2193 => (x"13",x"4b",x"71",x"1e"),
  2194 => (x"cb",x"02",x"9a",x"4a"),
  2195 => (x"fe",x"49",x"72",x"87"),
  2196 => (x"4a",x"13",x"87",x"e7"),
  2197 => (x"87",x"f5",x"05",x"9a"),
  2198 => (x"1e",x"87",x"da",x"fe"),
  2199 => (x"bf",x"ee",x"d9",x"c4"),
  2200 => (x"ee",x"d9",x"c4",x"49"),
  2201 => (x"78",x"a1",x"c1",x"48"),
  2202 => (x"a9",x"b7",x"c0",x"c4"),
  2203 => (x"ff",x"87",x"db",x"03"),
  2204 => (x"d9",x"c4",x"48",x"d4"),
  2205 => (x"c4",x"78",x"bf",x"f2"),
  2206 => (x"49",x"bf",x"ee",x"d9"),
  2207 => (x"48",x"ee",x"d9",x"c4"),
  2208 => (x"c4",x"78",x"a1",x"c1"),
  2209 => (x"04",x"a9",x"b7",x"c0"),
  2210 => (x"d0",x"ff",x"87",x"e5"),
  2211 => (x"c4",x"78",x"c8",x"48"),
  2212 => (x"c0",x"48",x"fa",x"d9"),
  2213 => (x"00",x"4f",x"26",x"78"),
  2214 => (x"00",x"00",x"00",x"00"),
  2215 => (x"00",x"00",x"00",x"00"),
  2216 => (x"5f",x"5f",x"00",x"00"),
  2217 => (x"00",x"00",x"00",x"00"),
  2218 => (x"03",x"00",x"03",x"03"),
  2219 => (x"14",x"00",x"00",x"03"),
  2220 => (x"7f",x"14",x"7f",x"7f"),
  2221 => (x"00",x"00",x"14",x"7f"),
  2222 => (x"6b",x"6b",x"2e",x"24"),
  2223 => (x"4c",x"00",x"12",x"3a"),
  2224 => (x"6c",x"18",x"36",x"6a"),
  2225 => (x"30",x"00",x"32",x"56"),
  2226 => (x"77",x"59",x"4f",x"7e"),
  2227 => (x"00",x"40",x"68",x"3a"),
  2228 => (x"03",x"07",x"04",x"00"),
  2229 => (x"00",x"00",x"00",x"00"),
  2230 => (x"63",x"3e",x"1c",x"00"),
  2231 => (x"00",x"00",x"00",x"41"),
  2232 => (x"3e",x"63",x"41",x"00"),
  2233 => (x"08",x"00",x"00",x"1c"),
  2234 => (x"1c",x"1c",x"3e",x"2a"),
  2235 => (x"00",x"08",x"2a",x"3e"),
  2236 => (x"3e",x"3e",x"08",x"08"),
  2237 => (x"00",x"00",x"08",x"08"),
  2238 => (x"60",x"e0",x"80",x"00"),
  2239 => (x"00",x"00",x"00",x"00"),
  2240 => (x"08",x"08",x"08",x"08"),
  2241 => (x"00",x"00",x"08",x"08"),
  2242 => (x"60",x"60",x"00",x"00"),
  2243 => (x"40",x"00",x"00",x"00"),
  2244 => (x"0c",x"18",x"30",x"60"),
  2245 => (x"00",x"01",x"03",x"06"),
  2246 => (x"4d",x"59",x"7f",x"3e"),
  2247 => (x"00",x"00",x"3e",x"7f"),
  2248 => (x"7f",x"7f",x"06",x"04"),
  2249 => (x"00",x"00",x"00",x"00"),
  2250 => (x"59",x"71",x"63",x"42"),
  2251 => (x"00",x"00",x"46",x"4f"),
  2252 => (x"49",x"49",x"63",x"22"),
  2253 => (x"18",x"00",x"36",x"7f"),
  2254 => (x"7f",x"13",x"16",x"1c"),
  2255 => (x"00",x"00",x"10",x"7f"),
  2256 => (x"45",x"45",x"67",x"27"),
  2257 => (x"00",x"00",x"39",x"7d"),
  2258 => (x"49",x"4b",x"7e",x"3c"),
  2259 => (x"00",x"00",x"30",x"79"),
  2260 => (x"79",x"71",x"01",x"01"),
  2261 => (x"00",x"00",x"07",x"0f"),
  2262 => (x"49",x"49",x"7f",x"36"),
  2263 => (x"00",x"00",x"36",x"7f"),
  2264 => (x"69",x"49",x"4f",x"06"),
  2265 => (x"00",x"00",x"1e",x"3f"),
  2266 => (x"66",x"66",x"00",x"00"),
  2267 => (x"00",x"00",x"00",x"00"),
  2268 => (x"66",x"e6",x"80",x"00"),
  2269 => (x"00",x"00",x"00",x"00"),
  2270 => (x"14",x"14",x"08",x"08"),
  2271 => (x"00",x"00",x"22",x"22"),
  2272 => (x"14",x"14",x"14",x"14"),
  2273 => (x"00",x"00",x"14",x"14"),
  2274 => (x"14",x"14",x"22",x"22"),
  2275 => (x"00",x"00",x"08",x"08"),
  2276 => (x"59",x"51",x"03",x"02"),
  2277 => (x"3e",x"00",x"06",x"0f"),
  2278 => (x"55",x"5d",x"41",x"7f"),
  2279 => (x"00",x"00",x"1e",x"1f"),
  2280 => (x"09",x"09",x"7f",x"7e"),
  2281 => (x"00",x"00",x"7e",x"7f"),
  2282 => (x"49",x"49",x"7f",x"7f"),
  2283 => (x"00",x"00",x"36",x"7f"),
  2284 => (x"41",x"63",x"3e",x"1c"),
  2285 => (x"00",x"00",x"41",x"41"),
  2286 => (x"63",x"41",x"7f",x"7f"),
  2287 => (x"00",x"00",x"1c",x"3e"),
  2288 => (x"49",x"49",x"7f",x"7f"),
  2289 => (x"00",x"00",x"41",x"41"),
  2290 => (x"09",x"09",x"7f",x"7f"),
  2291 => (x"00",x"00",x"01",x"01"),
  2292 => (x"49",x"41",x"7f",x"3e"),
  2293 => (x"00",x"00",x"7a",x"7b"),
  2294 => (x"08",x"08",x"7f",x"7f"),
  2295 => (x"00",x"00",x"7f",x"7f"),
  2296 => (x"7f",x"7f",x"41",x"00"),
  2297 => (x"00",x"00",x"00",x"41"),
  2298 => (x"40",x"40",x"60",x"20"),
  2299 => (x"7f",x"00",x"3f",x"7f"),
  2300 => (x"36",x"1c",x"08",x"7f"),
  2301 => (x"00",x"00",x"41",x"63"),
  2302 => (x"40",x"40",x"7f",x"7f"),
  2303 => (x"7f",x"00",x"40",x"40"),
  2304 => (x"06",x"0c",x"06",x"7f"),
  2305 => (x"7f",x"00",x"7f",x"7f"),
  2306 => (x"18",x"0c",x"06",x"7f"),
  2307 => (x"00",x"00",x"7f",x"7f"),
  2308 => (x"41",x"41",x"7f",x"3e"),
  2309 => (x"00",x"00",x"3e",x"7f"),
  2310 => (x"09",x"09",x"7f",x"7f"),
  2311 => (x"3e",x"00",x"06",x"0f"),
  2312 => (x"7f",x"61",x"41",x"7f"),
  2313 => (x"00",x"00",x"40",x"7e"),
  2314 => (x"19",x"09",x"7f",x"7f"),
  2315 => (x"00",x"00",x"66",x"7f"),
  2316 => (x"59",x"4d",x"6f",x"26"),
  2317 => (x"00",x"00",x"32",x"7b"),
  2318 => (x"7f",x"7f",x"01",x"01"),
  2319 => (x"00",x"00",x"01",x"01"),
  2320 => (x"40",x"40",x"7f",x"3f"),
  2321 => (x"00",x"00",x"3f",x"7f"),
  2322 => (x"70",x"70",x"3f",x"0f"),
  2323 => (x"7f",x"00",x"0f",x"3f"),
  2324 => (x"30",x"18",x"30",x"7f"),
  2325 => (x"41",x"00",x"7f",x"7f"),
  2326 => (x"1c",x"1c",x"36",x"63"),
  2327 => (x"01",x"41",x"63",x"36"),
  2328 => (x"7c",x"7c",x"06",x"03"),
  2329 => (x"61",x"01",x"03",x"06"),
  2330 => (x"47",x"4d",x"59",x"71"),
  2331 => (x"00",x"00",x"41",x"43"),
  2332 => (x"41",x"7f",x"7f",x"00"),
  2333 => (x"01",x"00",x"00",x"41"),
  2334 => (x"18",x"0c",x"06",x"03"),
  2335 => (x"00",x"40",x"60",x"30"),
  2336 => (x"7f",x"41",x"41",x"00"),
  2337 => (x"08",x"00",x"00",x"7f"),
  2338 => (x"06",x"03",x"06",x"0c"),
  2339 => (x"80",x"00",x"08",x"0c"),
  2340 => (x"80",x"80",x"80",x"80"),
  2341 => (x"00",x"00",x"80",x"80"),
  2342 => (x"07",x"03",x"00",x"00"),
  2343 => (x"00",x"00",x"00",x"04"),
  2344 => (x"54",x"54",x"74",x"20"),
  2345 => (x"00",x"00",x"78",x"7c"),
  2346 => (x"44",x"44",x"7f",x"7f"),
  2347 => (x"00",x"00",x"38",x"7c"),
  2348 => (x"44",x"44",x"7c",x"38"),
  2349 => (x"00",x"00",x"00",x"44"),
  2350 => (x"44",x"44",x"7c",x"38"),
  2351 => (x"00",x"00",x"7f",x"7f"),
  2352 => (x"54",x"54",x"7c",x"38"),
  2353 => (x"00",x"00",x"18",x"5c"),
  2354 => (x"05",x"7f",x"7e",x"04"),
  2355 => (x"00",x"00",x"00",x"05"),
  2356 => (x"a4",x"a4",x"bc",x"18"),
  2357 => (x"00",x"00",x"7c",x"fc"),
  2358 => (x"04",x"04",x"7f",x"7f"),
  2359 => (x"00",x"00",x"78",x"7c"),
  2360 => (x"7d",x"3d",x"00",x"00"),
  2361 => (x"00",x"00",x"00",x"40"),
  2362 => (x"fd",x"80",x"80",x"80"),
  2363 => (x"00",x"00",x"00",x"7d"),
  2364 => (x"38",x"10",x"7f",x"7f"),
  2365 => (x"00",x"00",x"44",x"6c"),
  2366 => (x"7f",x"3f",x"00",x"00"),
  2367 => (x"7c",x"00",x"00",x"40"),
  2368 => (x"0c",x"18",x"0c",x"7c"),
  2369 => (x"00",x"00",x"78",x"7c"),
  2370 => (x"04",x"04",x"7c",x"7c"),
  2371 => (x"00",x"00",x"78",x"7c"),
  2372 => (x"44",x"44",x"7c",x"38"),
  2373 => (x"00",x"00",x"38",x"7c"),
  2374 => (x"24",x"24",x"fc",x"fc"),
  2375 => (x"00",x"00",x"18",x"3c"),
  2376 => (x"24",x"24",x"3c",x"18"),
  2377 => (x"00",x"00",x"fc",x"fc"),
  2378 => (x"04",x"04",x"7c",x"7c"),
  2379 => (x"00",x"00",x"08",x"0c"),
  2380 => (x"54",x"54",x"5c",x"48"),
  2381 => (x"00",x"00",x"20",x"74"),
  2382 => (x"44",x"7f",x"3f",x"04"),
  2383 => (x"00",x"00",x"00",x"44"),
  2384 => (x"40",x"40",x"7c",x"3c"),
  2385 => (x"00",x"00",x"7c",x"7c"),
  2386 => (x"60",x"60",x"3c",x"1c"),
  2387 => (x"3c",x"00",x"1c",x"3c"),
  2388 => (x"60",x"30",x"60",x"7c"),
  2389 => (x"44",x"00",x"3c",x"7c"),
  2390 => (x"38",x"10",x"38",x"6c"),
  2391 => (x"00",x"00",x"44",x"6c"),
  2392 => (x"60",x"e0",x"bc",x"1c"),
  2393 => (x"00",x"00",x"1c",x"3c"),
  2394 => (x"5c",x"74",x"64",x"44"),
  2395 => (x"00",x"00",x"44",x"4c"),
  2396 => (x"77",x"3e",x"08",x"08"),
  2397 => (x"00",x"00",x"41",x"41"),
  2398 => (x"7f",x"7f",x"00",x"00"),
  2399 => (x"00",x"00",x"00",x"00"),
  2400 => (x"3e",x"77",x"41",x"41"),
  2401 => (x"02",x"00",x"08",x"08"),
  2402 => (x"02",x"03",x"01",x"01"),
  2403 => (x"7f",x"00",x"01",x"02"),
  2404 => (x"7f",x"7f",x"7f",x"7f"),
  2405 => (x"08",x"00",x"7f",x"7f"),
  2406 => (x"3e",x"1c",x"1c",x"08"),
  2407 => (x"7f",x"7f",x"7f",x"3e"),
  2408 => (x"1c",x"3e",x"3e",x"7f"),
  2409 => (x"00",x"08",x"08",x"1c"),
  2410 => (x"7c",x"7c",x"18",x"10"),
  2411 => (x"00",x"00",x"10",x"18"),
  2412 => (x"7c",x"7c",x"30",x"10"),
  2413 => (x"10",x"00",x"10",x"30"),
  2414 => (x"78",x"60",x"60",x"30"),
  2415 => (x"42",x"00",x"06",x"1e"),
  2416 => (x"3c",x"18",x"3c",x"66"),
  2417 => (x"78",x"00",x"42",x"66"),
  2418 => (x"c6",x"c2",x"6a",x"38"),
  2419 => (x"60",x"00",x"38",x"6c"),
  2420 => (x"00",x"60",x"00",x"00"),
  2421 => (x"0e",x"00",x"60",x"00"),
  2422 => (x"5d",x"5c",x"5b",x"5e"),
  2423 => (x"4c",x"71",x"1e",x"0e"),
  2424 => (x"bf",x"cb",x"da",x"c4"),
  2425 => (x"c0",x"4b",x"c0",x"4d"),
  2426 => (x"02",x"ab",x"74",x"1e"),
  2427 => (x"a6",x"c4",x"87",x"c7"),
  2428 => (x"c5",x"78",x"c0",x"48"),
  2429 => (x"48",x"a6",x"c4",x"87"),
  2430 => (x"66",x"c4",x"78",x"c1"),
  2431 => (x"ee",x"49",x"73",x"1e"),
  2432 => (x"86",x"c8",x"87",x"df"),
  2433 => (x"ef",x"49",x"e0",x"c0"),
  2434 => (x"a5",x"c4",x"87",x"ef"),
  2435 => (x"f0",x"49",x"6a",x"4a"),
  2436 => (x"c6",x"f1",x"87",x"f0"),
  2437 => (x"c1",x"85",x"cb",x"87"),
  2438 => (x"ab",x"b7",x"c8",x"83"),
  2439 => (x"87",x"c7",x"ff",x"04"),
  2440 => (x"26",x"4d",x"26",x"26"),
  2441 => (x"26",x"4b",x"26",x"4c"),
  2442 => (x"4a",x"71",x"1e",x"4f"),
  2443 => (x"5a",x"cf",x"da",x"c4"),
  2444 => (x"48",x"cf",x"da",x"c4"),
  2445 => (x"fe",x"49",x"78",x"c7"),
  2446 => (x"4f",x"26",x"87",x"dd"),
  2447 => (x"71",x"1e",x"73",x"1e"),
  2448 => (x"aa",x"b7",x"c0",x"4a"),
  2449 => (x"c2",x"87",x"d3",x"03"),
  2450 => (x"05",x"bf",x"e5",x"e6"),
  2451 => (x"4b",x"c1",x"87",x"c4"),
  2452 => (x"4b",x"c0",x"87",x"c2"),
  2453 => (x"5b",x"e9",x"e6",x"c2"),
  2454 => (x"e6",x"c2",x"87",x"c4"),
  2455 => (x"e6",x"c2",x"5a",x"e9"),
  2456 => (x"c1",x"4a",x"bf",x"e5"),
  2457 => (x"a2",x"c0",x"c1",x"9a"),
  2458 => (x"87",x"e8",x"ec",x"49"),
  2459 => (x"e6",x"c2",x"48",x"fc"),
  2460 => (x"fe",x"78",x"bf",x"e5"),
  2461 => (x"c2",x"1e",x"87",x"ef"),
  2462 => (x"48",x"bf",x"e5",x"e6"),
  2463 => (x"71",x"1e",x"4f",x"26"),
  2464 => (x"1e",x"66",x"c4",x"4a"),
  2465 => (x"f9",x"e9",x"49",x"72"),
  2466 => (x"4f",x"26",x"26",x"87"),
  2467 => (x"e5",x"e6",x"c2",x"1e"),
  2468 => (x"d8",x"c1",x"49",x"bf"),
  2469 => (x"da",x"c4",x"87",x"c5"),
  2470 => (x"bf",x"e8",x"48",x"c3"),
  2471 => (x"ff",x"d9",x"c4",x"78"),
  2472 => (x"78",x"bf",x"ec",x"48"),
  2473 => (x"bf",x"c3",x"da",x"c4"),
  2474 => (x"ff",x"c3",x"49",x"4a"),
  2475 => (x"2a",x"b7",x"c8",x"99"),
  2476 => (x"b0",x"71",x"48",x"72"),
  2477 => (x"58",x"cb",x"da",x"c4"),
  2478 => (x"5e",x"0e",x"4f",x"26"),
  2479 => (x"0e",x"5d",x"5c",x"5b"),
  2480 => (x"c7",x"ff",x"4b",x"71"),
  2481 => (x"fe",x"d9",x"c4",x"87"),
  2482 => (x"73",x"50",x"c0",x"48"),
  2483 => (x"fe",x"de",x"ff",x"49"),
  2484 => (x"4c",x"49",x"70",x"87"),
  2485 => (x"ee",x"cb",x"9c",x"c2"),
  2486 => (x"87",x"d1",x"cb",x"49"),
  2487 => (x"c4",x"4d",x"49",x"70"),
  2488 => (x"bf",x"97",x"fe",x"d9"),
  2489 => (x"87",x"e4",x"c1",x"05"),
  2490 => (x"c4",x"49",x"66",x"d0"),
  2491 => (x"99",x"bf",x"c7",x"da"),
  2492 => (x"d4",x"87",x"d7",x"05"),
  2493 => (x"d9",x"c4",x"49",x"66"),
  2494 => (x"05",x"99",x"bf",x"ff"),
  2495 => (x"49",x"73",x"87",x"cc"),
  2496 => (x"87",x"cb",x"de",x"ff"),
  2497 => (x"c1",x"02",x"98",x"70"),
  2498 => (x"4c",x"c1",x"87",x"c2"),
  2499 => (x"75",x"87",x"fd",x"fd"),
  2500 => (x"87",x"e5",x"ca",x"49"),
  2501 => (x"c6",x"02",x"98",x"70"),
  2502 => (x"fe",x"d9",x"c4",x"87"),
  2503 => (x"c4",x"50",x"c1",x"48"),
  2504 => (x"bf",x"97",x"fe",x"d9"),
  2505 => (x"87",x"e4",x"c0",x"05"),
  2506 => (x"bf",x"c7",x"da",x"c4"),
  2507 => (x"99",x"66",x"d0",x"49"),
  2508 => (x"87",x"d6",x"ff",x"05"),
  2509 => (x"bf",x"ff",x"d9",x"c4"),
  2510 => (x"99",x"66",x"d4",x"49"),
  2511 => (x"87",x"ca",x"ff",x"05"),
  2512 => (x"dd",x"ff",x"49",x"73"),
  2513 => (x"98",x"70",x"87",x"c9"),
  2514 => (x"87",x"fe",x"fe",x"05"),
  2515 => (x"d0",x"fb",x"48",x"74"),
  2516 => (x"5b",x"5e",x"0e",x"87"),
  2517 => (x"f4",x"0e",x"5d",x"5c"),
  2518 => (x"4c",x"4d",x"c0",x"86"),
  2519 => (x"c4",x"7e",x"bf",x"ec"),
  2520 => (x"da",x"c4",x"48",x"a6"),
  2521 => (x"c1",x"78",x"bf",x"cb"),
  2522 => (x"c3",x"1e",x"c0",x"1e"),
  2523 => (x"c9",x"fd",x"49",x"fc"),
  2524 => (x"70",x"86",x"c8",x"87"),
  2525 => (x"87",x"ce",x"02",x"98"),
  2526 => (x"ff",x"fa",x"49",x"ff"),
  2527 => (x"49",x"da",x"c1",x"87"),
  2528 => (x"87",x"cb",x"dc",x"ff"),
  2529 => (x"d9",x"c4",x"4d",x"c1"),
  2530 => (x"02",x"bf",x"97",x"fe"),
  2531 => (x"f8",x"c0",x"87",x"c4"),
  2532 => (x"da",x"c4",x"87",x"ef"),
  2533 => (x"c2",x"4b",x"bf",x"c3"),
  2534 => (x"05",x"bf",x"e5",x"e6"),
  2535 => (x"c3",x"87",x"eb",x"c0"),
  2536 => (x"db",x"ff",x"49",x"fd"),
  2537 => (x"fa",x"c3",x"87",x"e9"),
  2538 => (x"e2",x"db",x"ff",x"49"),
  2539 => (x"c3",x"49",x"73",x"87"),
  2540 => (x"1e",x"71",x"99",x"ff"),
  2541 => (x"c5",x"fb",x"49",x"c0"),
  2542 => (x"c8",x"49",x"73",x"87"),
  2543 => (x"1e",x"71",x"29",x"b7"),
  2544 => (x"f9",x"fa",x"49",x"c1"),
  2545 => (x"c6",x"86",x"c8",x"87"),
  2546 => (x"da",x"c4",x"87",x"c1"),
  2547 => (x"9b",x"4b",x"bf",x"c7"),
  2548 => (x"c2",x"87",x"dd",x"02"),
  2549 => (x"49",x"bf",x"e1",x"e6"),
  2550 => (x"70",x"87",x"de",x"c7"),
  2551 => (x"87",x"c4",x"05",x"98"),
  2552 => (x"87",x"d2",x"4b",x"c0"),
  2553 => (x"c7",x"49",x"e0",x"c2"),
  2554 => (x"e6",x"c2",x"87",x"c3"),
  2555 => (x"87",x"c6",x"58",x"e5"),
  2556 => (x"48",x"e1",x"e6",x"c2"),
  2557 => (x"49",x"73",x"78",x"c0"),
  2558 => (x"ce",x"05",x"99",x"c2"),
  2559 => (x"49",x"eb",x"c3",x"87"),
  2560 => (x"87",x"cb",x"da",x"ff"),
  2561 => (x"99",x"c2",x"49",x"70"),
  2562 => (x"fb",x"87",x"c2",x"02"),
  2563 => (x"c1",x"49",x"73",x"4c"),
  2564 => (x"87",x"ce",x"05",x"99"),
  2565 => (x"ff",x"49",x"f4",x"c3"),
  2566 => (x"70",x"87",x"f4",x"d9"),
  2567 => (x"02",x"99",x"c2",x"49"),
  2568 => (x"4c",x"fa",x"87",x"c2"),
  2569 => (x"99",x"c8",x"49",x"73"),
  2570 => (x"c3",x"87",x"ce",x"05"),
  2571 => (x"d9",x"ff",x"49",x"f5"),
  2572 => (x"49",x"70",x"87",x"dd"),
  2573 => (x"d5",x"02",x"99",x"c2"),
  2574 => (x"cf",x"da",x"c4",x"87"),
  2575 => (x"87",x"ca",x"02",x"bf"),
  2576 => (x"c4",x"88",x"c1",x"48"),
  2577 => (x"c0",x"58",x"d3",x"da"),
  2578 => (x"4c",x"ff",x"87",x"c2"),
  2579 => (x"49",x"73",x"4d",x"c1"),
  2580 => (x"ce",x"05",x"99",x"c4"),
  2581 => (x"49",x"f2",x"c3",x"87"),
  2582 => (x"87",x"f3",x"d8",x"ff"),
  2583 => (x"99",x"c2",x"49",x"70"),
  2584 => (x"c4",x"87",x"dc",x"02"),
  2585 => (x"7e",x"bf",x"cf",x"da"),
  2586 => (x"a8",x"b7",x"c7",x"48"),
  2587 => (x"87",x"cb",x"c0",x"03"),
  2588 => (x"80",x"c1",x"48",x"6e"),
  2589 => (x"58",x"d3",x"da",x"c4"),
  2590 => (x"fe",x"87",x"c2",x"c0"),
  2591 => (x"c3",x"4d",x"c1",x"4c"),
  2592 => (x"d8",x"ff",x"49",x"fd"),
  2593 => (x"49",x"70",x"87",x"c9"),
  2594 => (x"c0",x"02",x"99",x"c2"),
  2595 => (x"da",x"c4",x"87",x"d5"),
  2596 => (x"c0",x"02",x"bf",x"cf"),
  2597 => (x"da",x"c4",x"87",x"c9"),
  2598 => (x"78",x"c0",x"48",x"cf"),
  2599 => (x"fd",x"87",x"c2",x"c0"),
  2600 => (x"c3",x"4d",x"c1",x"4c"),
  2601 => (x"d7",x"ff",x"49",x"fa"),
  2602 => (x"49",x"70",x"87",x"e5"),
  2603 => (x"c0",x"02",x"99",x"c2"),
  2604 => (x"da",x"c4",x"87",x"d9"),
  2605 => (x"c7",x"48",x"bf",x"cf"),
  2606 => (x"c0",x"03",x"a8",x"b7"),
  2607 => (x"da",x"c4",x"87",x"c9"),
  2608 => (x"78",x"c7",x"48",x"cf"),
  2609 => (x"fc",x"87",x"c2",x"c0"),
  2610 => (x"c0",x"4d",x"c1",x"4c"),
  2611 => (x"c0",x"03",x"ac",x"b7"),
  2612 => (x"66",x"c4",x"87",x"d1"),
  2613 => (x"82",x"d8",x"c1",x"4a"),
  2614 => (x"c6",x"c0",x"02",x"6a"),
  2615 => (x"74",x"4b",x"6a",x"87"),
  2616 => (x"c0",x"0f",x"73",x"49"),
  2617 => (x"1e",x"f0",x"c3",x"1e"),
  2618 => (x"f7",x"49",x"da",x"c1"),
  2619 => (x"86",x"c8",x"87",x"cc"),
  2620 => (x"c0",x"02",x"98",x"70"),
  2621 => (x"a6",x"c8",x"87",x"e2"),
  2622 => (x"cf",x"da",x"c4",x"48"),
  2623 => (x"66",x"c8",x"78",x"bf"),
  2624 => (x"c4",x"91",x"cb",x"49"),
  2625 => (x"80",x"71",x"48",x"66"),
  2626 => (x"bf",x"6e",x"7e",x"70"),
  2627 => (x"87",x"c8",x"c0",x"02"),
  2628 => (x"c8",x"4b",x"bf",x"6e"),
  2629 => (x"0f",x"73",x"49",x"66"),
  2630 => (x"c0",x"02",x"9d",x"75"),
  2631 => (x"da",x"c4",x"87",x"c8"),
  2632 => (x"f2",x"49",x"bf",x"cf"),
  2633 => (x"e6",x"c2",x"87",x"f1"),
  2634 => (x"c0",x"02",x"bf",x"e9"),
  2635 => (x"c2",x"49",x"87",x"dd"),
  2636 => (x"98",x"70",x"87",x"c7"),
  2637 => (x"87",x"d3",x"c0",x"02"),
  2638 => (x"bf",x"cf",x"da",x"c4"),
  2639 => (x"87",x"d7",x"f2",x"49"),
  2640 => (x"f7",x"f3",x"49",x"c0"),
  2641 => (x"e9",x"e6",x"c2",x"87"),
  2642 => (x"f4",x"78",x"c0",x"48"),
  2643 => (x"87",x"d1",x"f3",x"8e"),
  2644 => (x"5c",x"5b",x"5e",x"0e"),
  2645 => (x"71",x"1e",x"0e",x"5d"),
  2646 => (x"cb",x"da",x"c4",x"4c"),
  2647 => (x"cd",x"c1",x"49",x"bf"),
  2648 => (x"d1",x"c1",x"4d",x"a1"),
  2649 => (x"74",x"7e",x"69",x"81"),
  2650 => (x"87",x"cf",x"02",x"9c"),
  2651 => (x"74",x"4b",x"a5",x"c4"),
  2652 => (x"cb",x"da",x"c4",x"7b"),
  2653 => (x"f0",x"f2",x"49",x"bf"),
  2654 => (x"74",x"7b",x"6e",x"87"),
  2655 => (x"87",x"c4",x"05",x"9c"),
  2656 => (x"87",x"c2",x"4b",x"c0"),
  2657 => (x"49",x"73",x"4b",x"c1"),
  2658 => (x"d4",x"87",x"f1",x"f2"),
  2659 => (x"87",x"c7",x"02",x"66"),
  2660 => (x"70",x"87",x"da",x"49"),
  2661 => (x"c0",x"87",x"c2",x"4a"),
  2662 => (x"ed",x"e6",x"c2",x"4a"),
  2663 => (x"c0",x"f2",x"26",x"5a"),
  2664 => (x"00",x"00",x"00",x"87"),
  2665 => (x"00",x"00",x"00",x"00"),
  2666 => (x"00",x"00",x"00",x"00"),
  2667 => (x"4a",x"71",x"1e",x"00"),
  2668 => (x"49",x"bf",x"c8",x"ff"),
  2669 => (x"26",x"48",x"a1",x"72"),
  2670 => (x"c8",x"ff",x"1e",x"4f"),
  2671 => (x"c0",x"fe",x"89",x"bf"),
  2672 => (x"c0",x"c0",x"c0",x"c0"),
  2673 => (x"87",x"c4",x"01",x"a9"),
  2674 => (x"87",x"c2",x"4a",x"c0"),
  2675 => (x"48",x"72",x"4a",x"c1"),
  2676 => (x"5e",x"0e",x"4f",x"26"),
  2677 => (x"0e",x"5d",x"5c",x"5b"),
  2678 => (x"d4",x"ff",x"4b",x"71"),
  2679 => (x"48",x"66",x"d0",x"4c"),
  2680 => (x"49",x"d6",x"78",x"c0"),
  2681 => (x"87",x"e0",x"db",x"ff"),
  2682 => (x"6c",x"7c",x"ff",x"c3"),
  2683 => (x"99",x"ff",x"c3",x"49"),
  2684 => (x"c3",x"49",x"4d",x"71"),
  2685 => (x"e0",x"c1",x"99",x"f0"),
  2686 => (x"87",x"cb",x"05",x"a9"),
  2687 => (x"6c",x"7c",x"ff",x"c3"),
  2688 => (x"d0",x"98",x"c3",x"48"),
  2689 => (x"c3",x"78",x"08",x"66"),
  2690 => (x"4a",x"6c",x"7c",x"ff"),
  2691 => (x"c3",x"31",x"c8",x"49"),
  2692 => (x"4a",x"6c",x"7c",x"ff"),
  2693 => (x"49",x"72",x"b2",x"71"),
  2694 => (x"ff",x"c3",x"31",x"c8"),
  2695 => (x"71",x"4a",x"6c",x"7c"),
  2696 => (x"c8",x"49",x"72",x"b2"),
  2697 => (x"7c",x"ff",x"c3",x"31"),
  2698 => (x"b2",x"71",x"4a",x"6c"),
  2699 => (x"c0",x"48",x"d0",x"ff"),
  2700 => (x"9b",x"73",x"78",x"e0"),
  2701 => (x"72",x"87",x"c2",x"02"),
  2702 => (x"26",x"48",x"75",x"7b"),
  2703 => (x"26",x"4c",x"26",x"4d"),
  2704 => (x"1e",x"4f",x"26",x"4b"),
  2705 => (x"5e",x"0e",x"4f",x"26"),
  2706 => (x"f8",x"0e",x"5c",x"5b"),
  2707 => (x"c8",x"1e",x"76",x"86"),
  2708 => (x"fd",x"fd",x"49",x"a6"),
  2709 => (x"70",x"86",x"c4",x"87"),
  2710 => (x"c2",x"48",x"6e",x"4b"),
  2711 => (x"f4",x"c2",x"03",x"a8"),
  2712 => (x"c3",x"4a",x"73",x"87"),
  2713 => (x"d0",x"c1",x"9a",x"f0"),
  2714 => (x"87",x"c7",x"02",x"aa"),
  2715 => (x"05",x"aa",x"e0",x"c1"),
  2716 => (x"73",x"87",x"e2",x"c2"),
  2717 => (x"02",x"99",x"c8",x"49"),
  2718 => (x"c6",x"ff",x"87",x"c3"),
  2719 => (x"c3",x"4c",x"73",x"87"),
  2720 => (x"05",x"ac",x"c2",x"9c"),
  2721 => (x"c4",x"87",x"c4",x"c1"),
  2722 => (x"31",x"c9",x"49",x"66"),
  2723 => (x"66",x"c4",x"1e",x"71"),
  2724 => (x"92",x"c8",x"c1",x"4a"),
  2725 => (x"49",x"d3",x"da",x"c4"),
  2726 => (x"c2",x"fe",x"81",x"72"),
  2727 => (x"49",x"d8",x"87",x"d6"),
  2728 => (x"87",x"e4",x"d8",x"ff"),
  2729 => (x"c4",x"1e",x"c0",x"c8"),
  2730 => (x"fd",x"49",x"da",x"c7"),
  2731 => (x"ff",x"87",x"e2",x"da"),
  2732 => (x"e0",x"c0",x"48",x"d0"),
  2733 => (x"da",x"c7",x"c4",x"78"),
  2734 => (x"4a",x"66",x"cc",x"1e"),
  2735 => (x"c4",x"92",x"c8",x"c1"),
  2736 => (x"72",x"49",x"d3",x"da"),
  2737 => (x"e0",x"fd",x"fd",x"81"),
  2738 => (x"c1",x"86",x"cc",x"87"),
  2739 => (x"c4",x"c1",x"05",x"ac"),
  2740 => (x"49",x"66",x"c4",x"87"),
  2741 => (x"1e",x"71",x"31",x"c9"),
  2742 => (x"c1",x"4a",x"66",x"c4"),
  2743 => (x"da",x"c4",x"92",x"c8"),
  2744 => (x"81",x"72",x"49",x"d3"),
  2745 => (x"87",x"cc",x"c1",x"fe"),
  2746 => (x"1e",x"da",x"c7",x"c4"),
  2747 => (x"c1",x"4a",x"66",x"c8"),
  2748 => (x"da",x"c4",x"92",x"c8"),
  2749 => (x"81",x"72",x"49",x"d3"),
  2750 => (x"87",x"de",x"fb",x"fd"),
  2751 => (x"d7",x"ff",x"49",x"d7"),
  2752 => (x"c0",x"c8",x"87",x"c6"),
  2753 => (x"da",x"c7",x"c4",x"1e"),
  2754 => (x"dd",x"d8",x"fd",x"49"),
  2755 => (x"ff",x"86",x"cc",x"87"),
  2756 => (x"e0",x"c0",x"48",x"d0"),
  2757 => (x"fc",x"8e",x"f8",x"78"),
  2758 => (x"5e",x"0e",x"87",x"e3"),
  2759 => (x"0e",x"5d",x"5c",x"5b"),
  2760 => (x"ff",x"4d",x"71",x"1e"),
  2761 => (x"66",x"d4",x"4c",x"d4"),
  2762 => (x"b7",x"c3",x"48",x"7e"),
  2763 => (x"87",x"c5",x"06",x"a8"),
  2764 => (x"e3",x"c1",x"48",x"c0"),
  2765 => (x"fe",x"49",x"75",x"87"),
  2766 => (x"75",x"87",x"e6",x"d0"),
  2767 => (x"4b",x"66",x"c4",x"1e"),
  2768 => (x"c4",x"93",x"c8",x"c1"),
  2769 => (x"73",x"83",x"d3",x"da"),
  2770 => (x"e6",x"f4",x"fd",x"49"),
  2771 => (x"6b",x"83",x"c8",x"87"),
  2772 => (x"48",x"d0",x"ff",x"4b"),
  2773 => (x"dd",x"78",x"e1",x"c8"),
  2774 => (x"c3",x"49",x"73",x"7c"),
  2775 => (x"7c",x"71",x"99",x"ff"),
  2776 => (x"b7",x"c8",x"49",x"73"),
  2777 => (x"99",x"ff",x"c3",x"29"),
  2778 => (x"49",x"73",x"7c",x"71"),
  2779 => (x"c3",x"29",x"b7",x"d0"),
  2780 => (x"7c",x"71",x"99",x"ff"),
  2781 => (x"b7",x"d8",x"49",x"73"),
  2782 => (x"c0",x"7c",x"71",x"29"),
  2783 => (x"7c",x"7c",x"7c",x"7c"),
  2784 => (x"7c",x"7c",x"7c",x"7c"),
  2785 => (x"7c",x"7c",x"7c",x"7c"),
  2786 => (x"c4",x"78",x"e0",x"c0"),
  2787 => (x"49",x"dc",x"1e",x"66"),
  2788 => (x"87",x"d9",x"d5",x"ff"),
  2789 => (x"48",x"73",x"86",x"c8"),
  2790 => (x"87",x"df",x"fa",x"26"),
  2791 => (x"4a",x"d4",x"ff",x"1e"),
  2792 => (x"c8",x"48",x"d0",x"ff"),
  2793 => (x"f0",x"c3",x"78",x"c5"),
  2794 => (x"c0",x"7a",x"71",x"7a"),
  2795 => (x"7a",x"7a",x"7a",x"7a"),
  2796 => (x"4f",x"26",x"78",x"c4"),
  2797 => (x"4a",x"d4",x"ff",x"1e"),
  2798 => (x"c8",x"48",x"d0",x"ff"),
  2799 => (x"7a",x"c0",x"78",x"c5"),
  2800 => (x"7a",x"c0",x"49",x"6a"),
  2801 => (x"7a",x"7a",x"7a",x"7a"),
  2802 => (x"48",x"71",x"78",x"c4"),
  2803 => (x"73",x"1e",x"4f",x"26"),
  2804 => (x"c8",x"4b",x"71",x"1e"),
  2805 => (x"87",x"db",x"02",x"66"),
  2806 => (x"c1",x"4a",x"6b",x"97"),
  2807 => (x"69",x"97",x"49",x"a3"),
  2808 => (x"51",x"72",x"7b",x"97"),
  2809 => (x"c2",x"48",x"66",x"c8"),
  2810 => (x"58",x"a6",x"cc",x"88"),
  2811 => (x"98",x"70",x"83",x"c2"),
  2812 => (x"c4",x"87",x"e5",x"05"),
  2813 => (x"26",x"4d",x"26",x"87"),
  2814 => (x"26",x"4b",x"26",x"4c"),
  2815 => (x"5b",x"5e",x"0e",x"4f"),
  2816 => (x"e8",x"0e",x"5d",x"5c"),
  2817 => (x"59",x"a6",x"cc",x"86"),
  2818 => (x"4d",x"66",x"e8",x"c0"),
  2819 => (x"c4",x"95",x"dc",x"c1"),
  2820 => (x"c1",x"85",x"e3",x"dc"),
  2821 => (x"c4",x"7e",x"a5",x"c8"),
  2822 => (x"cc",x"c1",x"48",x"a6"),
  2823 => (x"66",x"c4",x"78",x"a5"),
  2824 => (x"bf",x"6e",x"4c",x"bf"),
  2825 => (x"85",x"d0",x"c1",x"94"),
  2826 => (x"66",x"c8",x"94",x"6d"),
  2827 => (x"c8",x"4a",x"c0",x"4b"),
  2828 => (x"d2",x"fd",x"49",x"c0"),
  2829 => (x"66",x"c8",x"87",x"c2"),
  2830 => (x"9f",x"c0",x"c1",x"48"),
  2831 => (x"49",x"66",x"c8",x"78"),
  2832 => (x"bf",x"6e",x"81",x"c2"),
  2833 => (x"66",x"c8",x"79",x"9f"),
  2834 => (x"c4",x"81",x"c6",x"49"),
  2835 => (x"79",x"9f",x"bf",x"66"),
  2836 => (x"cc",x"49",x"66",x"c8"),
  2837 => (x"79",x"9f",x"6d",x"81"),
  2838 => (x"d4",x"48",x"66",x"c8"),
  2839 => (x"58",x"a6",x"d0",x"80"),
  2840 => (x"48",x"e9",x"f4",x"c2"),
  2841 => (x"d4",x"49",x"66",x"cc"),
  2842 => (x"41",x"20",x"4a",x"a1"),
  2843 => (x"f9",x"05",x"aa",x"71"),
  2844 => (x"48",x"66",x"c8",x"87"),
  2845 => (x"d4",x"80",x"ee",x"c0"),
  2846 => (x"f4",x"c2",x"58",x"a6"),
  2847 => (x"66",x"d0",x"48",x"fe"),
  2848 => (x"4a",x"a1",x"c8",x"49"),
  2849 => (x"aa",x"71",x"41",x"20"),
  2850 => (x"c8",x"87",x"f9",x"05"),
  2851 => (x"f6",x"c0",x"48",x"66"),
  2852 => (x"58",x"a6",x"d8",x"80"),
  2853 => (x"48",x"c7",x"f5",x"c2"),
  2854 => (x"c0",x"49",x"66",x"d4"),
  2855 => (x"20",x"4a",x"a1",x"e8"),
  2856 => (x"05",x"aa",x"71",x"41"),
  2857 => (x"e8",x"c0",x"87",x"f9"),
  2858 => (x"49",x"66",x"d8",x"1e"),
  2859 => (x"cc",x"87",x"df",x"fc"),
  2860 => (x"de",x"c1",x"49",x"66"),
  2861 => (x"d0",x"c0",x"c8",x"81"),
  2862 => (x"66",x"cc",x"79",x"9f"),
  2863 => (x"81",x"e2",x"c1",x"49"),
  2864 => (x"79",x"9f",x"c0",x"c8"),
  2865 => (x"c1",x"49",x"66",x"cc"),
  2866 => (x"9f",x"c1",x"81",x"ea"),
  2867 => (x"49",x"66",x"cc",x"79"),
  2868 => (x"c4",x"81",x"ec",x"c1"),
  2869 => (x"79",x"9f",x"bf",x"66"),
  2870 => (x"c1",x"49",x"66",x"cc"),
  2871 => (x"66",x"c8",x"81",x"ee"),
  2872 => (x"cc",x"79",x"9f",x"bf"),
  2873 => (x"f0",x"c1",x"49",x"66"),
  2874 => (x"79",x"9f",x"6d",x"81"),
  2875 => (x"ff",x"cf",x"4b",x"74"),
  2876 => (x"4a",x"73",x"9b",x"ff"),
  2877 => (x"c1",x"49",x"66",x"cc"),
  2878 => (x"9f",x"72",x"81",x"f2"),
  2879 => (x"d0",x"4a",x"74",x"79"),
  2880 => (x"ff",x"ff",x"cf",x"2a"),
  2881 => (x"cc",x"4c",x"72",x"9a"),
  2882 => (x"f4",x"c1",x"49",x"66"),
  2883 => (x"79",x"9f",x"74",x"81"),
  2884 => (x"49",x"66",x"cc",x"73"),
  2885 => (x"73",x"81",x"f8",x"c1"),
  2886 => (x"cc",x"72",x"79",x"9f"),
  2887 => (x"fa",x"c1",x"49",x"66"),
  2888 => (x"79",x"9f",x"72",x"81"),
  2889 => (x"cc",x"fb",x"8e",x"e4"),
  2890 => (x"54",x"4d",x"69",x"87"),
  2891 => (x"69",x"4d",x"69",x"53"),
  2892 => (x"48",x"4d",x"69",x"6e"),
  2893 => (x"66",x"61",x"72",x"67"),
  2894 => (x"20",x"69",x"6c",x"64"),
  2895 => (x"31",x"2e",x"00",x"65"),
  2896 => (x"20",x"20",x"30",x"30"),
  2897 => (x"59",x"00",x"20",x"20"),
  2898 => (x"42",x"55",x"51",x"41"),
  2899 => (x"20",x"20",x"20",x"45"),
  2900 => (x"20",x"20",x"20",x"20"),
  2901 => (x"20",x"20",x"20",x"20"),
  2902 => (x"20",x"20",x"20",x"20"),
  2903 => (x"20",x"20",x"20",x"20"),
  2904 => (x"20",x"20",x"20",x"20"),
  2905 => (x"20",x"20",x"20",x"20"),
  2906 => (x"20",x"20",x"20",x"20"),
  2907 => (x"00",x"20",x"20",x"20"),
  2908 => (x"71",x"1e",x"73",x"1e"),
  2909 => (x"02",x"66",x"d4",x"4b"),
  2910 => (x"66",x"c8",x"87",x"d4"),
  2911 => (x"73",x"31",x"d8",x"49"),
  2912 => (x"72",x"32",x"c8",x"4a"),
  2913 => (x"66",x"cc",x"49",x"a1"),
  2914 => (x"c0",x"48",x"71",x"81"),
  2915 => (x"66",x"d0",x"87",x"e3"),
  2916 => (x"91",x"dc",x"c1",x"49"),
  2917 => (x"81",x"e3",x"dc",x"c4"),
  2918 => (x"4a",x"a1",x"cc",x"c1"),
  2919 => (x"92",x"73",x"4a",x"6a"),
  2920 => (x"c1",x"82",x"66",x"c8"),
  2921 => (x"49",x"69",x"81",x"d0"),
  2922 => (x"66",x"cc",x"91",x"72"),
  2923 => (x"71",x"89",x"c1",x"81"),
  2924 => (x"87",x"c5",x"f9",x"48"),
  2925 => (x"ff",x"4a",x"71",x"1e"),
  2926 => (x"d0",x"ff",x"49",x"d4"),
  2927 => (x"78",x"c5",x"c8",x"48"),
  2928 => (x"c0",x"79",x"d0",x"c2"),
  2929 => (x"79",x"79",x"79",x"79"),
  2930 => (x"79",x"79",x"79",x"79"),
  2931 => (x"79",x"c0",x"79",x"72"),
  2932 => (x"c0",x"79",x"66",x"c4"),
  2933 => (x"79",x"66",x"c8",x"79"),
  2934 => (x"66",x"cc",x"79",x"c0"),
  2935 => (x"d0",x"79",x"c0",x"79"),
  2936 => (x"79",x"c0",x"79",x"66"),
  2937 => (x"c4",x"79",x"66",x"d4"),
  2938 => (x"1e",x"4f",x"26",x"78"),
  2939 => (x"a2",x"c6",x"4a",x"71"),
  2940 => (x"49",x"69",x"97",x"49"),
  2941 => (x"71",x"99",x"f0",x"c3"),
  2942 => (x"1e",x"1e",x"c0",x"1e"),
  2943 => (x"1e",x"c0",x"1e",x"c1"),
  2944 => (x"87",x"f0",x"fe",x"49"),
  2945 => (x"f6",x"49",x"d0",x"c2"),
  2946 => (x"8e",x"ec",x"87",x"d2"),
  2947 => (x"c0",x"1e",x"4f",x"26"),
  2948 => (x"1e",x"1e",x"1e",x"1e"),
  2949 => (x"fe",x"49",x"c1",x"1e"),
  2950 => (x"d0",x"c2",x"87",x"da"),
  2951 => (x"87",x"fc",x"f5",x"49"),
  2952 => (x"4f",x"26",x"8e",x"ec"),
  2953 => (x"ff",x"4a",x"71",x"1e"),
  2954 => (x"c5",x"c8",x"48",x"d0"),
  2955 => (x"48",x"d4",x"ff",x"78"),
  2956 => (x"c0",x"78",x"e0",x"c2"),
  2957 => (x"78",x"78",x"78",x"78"),
  2958 => (x"1e",x"c0",x"c8",x"78"),
  2959 => (x"cb",x"fd",x"49",x"72"),
  2960 => (x"d0",x"ff",x"87",x"e8"),
  2961 => (x"26",x"78",x"c4",x"48"),
  2962 => (x"5e",x"0e",x"4f",x"26"),
  2963 => (x"0e",x"5d",x"5c",x"5b"),
  2964 => (x"4a",x"71",x"86",x"f8"),
  2965 => (x"c1",x"4b",x"a2",x"c2"),
  2966 => (x"a2",x"c3",x"7b",x"97"),
  2967 => (x"7c",x"97",x"c1",x"4c"),
  2968 => (x"51",x"c0",x"49",x"a2"),
  2969 => (x"c0",x"4d",x"a2",x"c4"),
  2970 => (x"a2",x"c5",x"7d",x"97"),
  2971 => (x"c0",x"48",x"6e",x"7e"),
  2972 => (x"48",x"a6",x"c4",x"50"),
  2973 => (x"c4",x"78",x"a2",x"c6"),
  2974 => (x"50",x"c0",x"48",x"66"),
  2975 => (x"c4",x"1e",x"66",x"d8"),
  2976 => (x"f5",x"49",x"da",x"c7"),
  2977 => (x"66",x"c8",x"87",x"f7"),
  2978 => (x"1e",x"49",x"bf",x"97"),
  2979 => (x"bf",x"97",x"66",x"c8"),
  2980 => (x"49",x"15",x"1e",x"49"),
  2981 => (x"1e",x"49",x"14",x"1e"),
  2982 => (x"c0",x"1e",x"49",x"13"),
  2983 => (x"87",x"d4",x"fc",x"49"),
  2984 => (x"f7",x"f3",x"49",x"c8"),
  2985 => (x"da",x"c7",x"c4",x"87"),
  2986 => (x"87",x"f8",x"fd",x"49"),
  2987 => (x"f3",x"49",x"d0",x"c2"),
  2988 => (x"8e",x"e0",x"87",x"ea"),
  2989 => (x"1e",x"87",x"fe",x"f4"),
  2990 => (x"a2",x"c6",x"4a",x"71"),
  2991 => (x"49",x"69",x"97",x"49"),
  2992 => (x"49",x"a2",x"c5",x"1e"),
  2993 => (x"1e",x"49",x"69",x"97"),
  2994 => (x"97",x"49",x"a2",x"c4"),
  2995 => (x"c3",x"1e",x"49",x"69"),
  2996 => (x"69",x"97",x"49",x"a2"),
  2997 => (x"a2",x"c2",x"1e",x"49"),
  2998 => (x"49",x"69",x"97",x"49"),
  2999 => (x"fb",x"49",x"c0",x"1e"),
  3000 => (x"d0",x"c2",x"87",x"d2"),
  3001 => (x"87",x"f4",x"f2",x"49"),
  3002 => (x"4f",x"26",x"8e",x"ec"),
  3003 => (x"71",x"1e",x"73",x"1e"),
  3004 => (x"4a",x"a3",x"c2",x"4b"),
  3005 => (x"c1",x"49",x"66",x"c8"),
  3006 => (x"dc",x"c4",x"91",x"dc"),
  3007 => (x"d4",x"c1",x"81",x"e3"),
  3008 => (x"c2",x"79",x"12",x"81"),
  3009 => (x"d3",x"f2",x"49",x"d0"),
  3010 => (x"87",x"ed",x"f3",x"87"),
  3011 => (x"71",x"1e",x"73",x"1e"),
  3012 => (x"49",x"a3",x"c6",x"4b"),
  3013 => (x"1e",x"49",x"69",x"97"),
  3014 => (x"97",x"49",x"a3",x"c5"),
  3015 => (x"c4",x"1e",x"49",x"69"),
  3016 => (x"69",x"97",x"49",x"a3"),
  3017 => (x"a3",x"c3",x"1e",x"49"),
  3018 => (x"49",x"69",x"97",x"49"),
  3019 => (x"49",x"a3",x"c2",x"1e"),
  3020 => (x"1e",x"49",x"69",x"97"),
  3021 => (x"12",x"4a",x"a3",x"c1"),
  3022 => (x"87",x"f8",x"f9",x"49"),
  3023 => (x"f1",x"49",x"d0",x"c2"),
  3024 => (x"8e",x"ec",x"87",x"da"),
  3025 => (x"0e",x"87",x"f2",x"f2"),
  3026 => (x"5d",x"5c",x"5b",x"5e"),
  3027 => (x"7e",x"71",x"1e",x"0e"),
  3028 => (x"81",x"c2",x"49",x"6e"),
  3029 => (x"6e",x"79",x"97",x"c1"),
  3030 => (x"c1",x"83",x"c3",x"4b"),
  3031 => (x"4a",x"6e",x"7b",x"97"),
  3032 => (x"97",x"c0",x"82",x"c1"),
  3033 => (x"c4",x"4c",x"6e",x"7a"),
  3034 => (x"7c",x"97",x"c0",x"84"),
  3035 => (x"85",x"c5",x"4d",x"6e"),
  3036 => (x"4d",x"6e",x"55",x"c0"),
  3037 => (x"6d",x"97",x"85",x"c6"),
  3038 => (x"1e",x"c0",x"1e",x"4d"),
  3039 => (x"1e",x"4c",x"6c",x"97"),
  3040 => (x"1e",x"4b",x"6b",x"97"),
  3041 => (x"1e",x"49",x"69",x"97"),
  3042 => (x"e7",x"f8",x"49",x"12"),
  3043 => (x"49",x"d0",x"c2",x"87"),
  3044 => (x"e8",x"87",x"c9",x"f0"),
  3045 => (x"87",x"dd",x"f1",x"8e"),
  3046 => (x"5c",x"5b",x"5e",x"0e"),
  3047 => (x"dc",x"ff",x"0e",x"5d"),
  3048 => (x"c3",x"4b",x"71",x"86"),
  3049 => (x"4c",x"11",x"49",x"a3"),
  3050 => (x"c5",x"4a",x"a3",x"c4"),
  3051 => (x"69",x"97",x"49",x"a3"),
  3052 => (x"97",x"31",x"c8",x"49"),
  3053 => (x"71",x"48",x"4a",x"6a"),
  3054 => (x"58",x"a6",x"d4",x"b0"),
  3055 => (x"6e",x"7e",x"a3",x"c6"),
  3056 => (x"4d",x"49",x"bf",x"97"),
  3057 => (x"48",x"71",x"9d",x"cf"),
  3058 => (x"d8",x"98",x"c0",x"c1"),
  3059 => (x"f0",x"48",x"58",x"a6"),
  3060 => (x"78",x"a3",x"c2",x"80"),
  3061 => (x"bf",x"97",x"66",x"c4"),
  3062 => (x"58",x"a6",x"d0",x"48"),
  3063 => (x"c0",x"1e",x"66",x"d4"),
  3064 => (x"74",x"1e",x"66",x"f8"),
  3065 => (x"c0",x"1e",x"75",x"1e"),
  3066 => (x"f6",x"49",x"66",x"e0"),
  3067 => (x"86",x"d0",x"87",x"c2"),
  3068 => (x"a6",x"dc",x"49",x"70"),
  3069 => (x"02",x"66",x"cc",x"59"),
  3070 => (x"c0",x"87",x"e4",x"c5"),
  3071 => (x"c5",x"02",x"66",x"f8"),
  3072 => (x"4a",x"66",x"cc",x"87"),
  3073 => (x"4a",x"c1",x"87",x"c2"),
  3074 => (x"f8",x"c0",x"4b",x"72"),
  3075 => (x"87",x"db",x"02",x"66"),
  3076 => (x"49",x"66",x"f4",x"c0"),
  3077 => (x"c4",x"91",x"dc",x"c1"),
  3078 => (x"c1",x"81",x"e3",x"dc"),
  3079 => (x"a6",x"c8",x"81",x"d4"),
  3080 => (x"c8",x"78",x"69",x"48"),
  3081 => (x"06",x"aa",x"b7",x"66"),
  3082 => (x"c8",x"4b",x"87",x"c1"),
  3083 => (x"87",x"ec",x"ed",x"49"),
  3084 => (x"70",x"87",x"c1",x"ee"),
  3085 => (x"05",x"99",x"c4",x"49"),
  3086 => (x"f7",x"ed",x"87",x"ca"),
  3087 => (x"c4",x"49",x"70",x"87"),
  3088 => (x"87",x"f6",x"02",x"99"),
  3089 => (x"88",x"c1",x"48",x"73"),
  3090 => (x"58",x"a6",x"e0",x"c0"),
  3091 => (x"dc",x"80",x"ec",x"48"),
  3092 => (x"9b",x"73",x"78",x"66"),
  3093 => (x"87",x"d0",x"c1",x"02"),
  3094 => (x"c1",x"48",x"66",x"cc"),
  3095 => (x"f0",x"c0",x"02",x"a8"),
  3096 => (x"66",x"f4",x"c0",x"87"),
  3097 => (x"91",x"dc",x"c1",x"49"),
  3098 => (x"4a",x"e3",x"dc",x"c4"),
  3099 => (x"d0",x"c1",x"82",x"71"),
  3100 => (x"ac",x"69",x"49",x"a2"),
  3101 => (x"c1",x"87",x"d8",x"05"),
  3102 => (x"cc",x"c1",x"85",x"4c"),
  3103 => (x"ad",x"69",x"49",x"a2"),
  3104 => (x"c0",x"87",x"ce",x"05"),
  3105 => (x"48",x"66",x"d0",x"4d"),
  3106 => (x"a6",x"d4",x"80",x"c1"),
  3107 => (x"c1",x"87",x"c2",x"58"),
  3108 => (x"48",x"66",x"cc",x"84"),
  3109 => (x"a6",x"d0",x"88",x"c1"),
  3110 => (x"49",x"66",x"c8",x"58"),
  3111 => (x"cc",x"88",x"c1",x"48"),
  3112 => (x"99",x"71",x"58",x"a6"),
  3113 => (x"87",x"f0",x"fe",x"05"),
  3114 => (x"d9",x"02",x"66",x"d4"),
  3115 => (x"d8",x"49",x"73",x"87"),
  3116 => (x"4a",x"71",x"81",x"66"),
  3117 => (x"72",x"9a",x"ff",x"c3"),
  3118 => (x"c8",x"4a",x"71",x"4c"),
  3119 => (x"a6",x"d4",x"2a",x"b7"),
  3120 => (x"29",x"b7",x"d8",x"5a"),
  3121 => (x"97",x"6e",x"4d",x"71"),
  3122 => (x"f0",x"c3",x"49",x"bf"),
  3123 => (x"71",x"b1",x"75",x"99"),
  3124 => (x"49",x"66",x"d4",x"1e"),
  3125 => (x"71",x"29",x"b7",x"c8"),
  3126 => (x"1e",x"66",x"d8",x"1e"),
  3127 => (x"66",x"d4",x"1e",x"74"),
  3128 => (x"1e",x"49",x"bf",x"97"),
  3129 => (x"cb",x"f3",x"49",x"c0"),
  3130 => (x"d0",x"86",x"d4",x"87"),
  3131 => (x"87",x"ec",x"ea",x"49"),
  3132 => (x"49",x"66",x"f4",x"c0"),
  3133 => (x"c4",x"91",x"dc",x"c1"),
  3134 => (x"71",x"48",x"e3",x"dc"),
  3135 => (x"58",x"a6",x"cc",x"80"),
  3136 => (x"c8",x"49",x"66",x"c8"),
  3137 => (x"c1",x"02",x"69",x"81"),
  3138 => (x"e0",x"c0",x"87",x"ca"),
  3139 => (x"66",x"dc",x"48",x"a6"),
  3140 => (x"02",x"9b",x"73",x"78"),
  3141 => (x"d8",x"87",x"c2",x"c1"),
  3142 => (x"31",x"c9",x"49",x"66"),
  3143 => (x"66",x"cc",x"1e",x"71"),
  3144 => (x"cf",x"e8",x"fd",x"49"),
  3145 => (x"d0",x"1e",x"c0",x"87"),
  3146 => (x"e2",x"fd",x"49",x"66"),
  3147 => (x"1e",x"c1",x"87",x"ec"),
  3148 => (x"fd",x"49",x"66",x"d4"),
  3149 => (x"cc",x"87",x"c9",x"e1"),
  3150 => (x"48",x"66",x"d8",x"86"),
  3151 => (x"a6",x"dc",x"80",x"c1"),
  3152 => (x"66",x"e0",x"c0",x"58"),
  3153 => (x"88",x"c1",x"48",x"49"),
  3154 => (x"58",x"a6",x"e4",x"c0"),
  3155 => (x"ff",x"05",x"99",x"71"),
  3156 => (x"87",x"c5",x"87",x"c5"),
  3157 => (x"c3",x"e9",x"49",x"c9"),
  3158 => (x"05",x"66",x"cc",x"87"),
  3159 => (x"c2",x"87",x"dc",x"fa"),
  3160 => (x"f7",x"e8",x"49",x"c0"),
  3161 => (x"8e",x"dc",x"ff",x"87"),
  3162 => (x"0e",x"87",x"ca",x"ea"),
  3163 => (x"5d",x"5c",x"5b",x"5e"),
  3164 => (x"71",x"86",x"e0",x"0e"),
  3165 => (x"49",x"a4",x"c3",x"4c"),
  3166 => (x"a6",x"d4",x"48",x"11"),
  3167 => (x"4a",x"a4",x"c4",x"58"),
  3168 => (x"97",x"49",x"a4",x"c5"),
  3169 => (x"31",x"c8",x"49",x"69"),
  3170 => (x"48",x"4a",x"6a",x"97"),
  3171 => (x"a6",x"d8",x"b0",x"71"),
  3172 => (x"7e",x"a4",x"c6",x"58"),
  3173 => (x"49",x"bf",x"97",x"6e"),
  3174 => (x"71",x"9d",x"cf",x"4d"),
  3175 => (x"98",x"c0",x"c1",x"48"),
  3176 => (x"48",x"58",x"a6",x"dc"),
  3177 => (x"a4",x"c2",x"80",x"ec"),
  3178 => (x"97",x"66",x"c4",x"78"),
  3179 => (x"66",x"d8",x"4b",x"bf"),
  3180 => (x"66",x"f4",x"c0",x"1e"),
  3181 => (x"1e",x"66",x"d8",x"1e"),
  3182 => (x"e4",x"c0",x"1e",x"75"),
  3183 => (x"ef",x"ee",x"49",x"66"),
  3184 => (x"70",x"86",x"d0",x"87"),
  3185 => (x"a6",x"e0",x"c0",x"49"),
  3186 => (x"05",x"9b",x"73",x"59"),
  3187 => (x"c0",x"c4",x"87",x"c3"),
  3188 => (x"e7",x"49",x"c4",x"4b"),
  3189 => (x"66",x"dc",x"87",x"c6"),
  3190 => (x"71",x"31",x"c9",x"49"),
  3191 => (x"66",x"f4",x"c0",x"1e"),
  3192 => (x"91",x"dc",x"c1",x"49"),
  3193 => (x"48",x"e3",x"dc",x"c4"),
  3194 => (x"a6",x"d4",x"80",x"71"),
  3195 => (x"49",x"66",x"d0",x"58"),
  3196 => (x"87",x"c0",x"e5",x"fd"),
  3197 => (x"9b",x"73",x"86",x"c4"),
  3198 => (x"87",x"df",x"c4",x"02"),
  3199 => (x"02",x"66",x"f4",x"c0"),
  3200 => (x"4a",x"73",x"87",x"c4"),
  3201 => (x"4a",x"c1",x"87",x"c2"),
  3202 => (x"f4",x"c0",x"4c",x"72"),
  3203 => (x"87",x"d3",x"02",x"66"),
  3204 => (x"c1",x"49",x"66",x"cc"),
  3205 => (x"a6",x"c8",x"81",x"d4"),
  3206 => (x"c8",x"78",x"69",x"48"),
  3207 => (x"06",x"aa",x"b7",x"66"),
  3208 => (x"74",x"4c",x"87",x"c1"),
  3209 => (x"d5",x"c2",x"02",x"9c"),
  3210 => (x"87",x"c8",x"e6",x"87"),
  3211 => (x"99",x"c8",x"49",x"70"),
  3212 => (x"e5",x"87",x"ca",x"05"),
  3213 => (x"49",x"70",x"87",x"fe"),
  3214 => (x"f6",x"02",x"99",x"c8"),
  3215 => (x"48",x"d0",x"ff",x"87"),
  3216 => (x"ff",x"78",x"c5",x"c8"),
  3217 => (x"f0",x"c2",x"48",x"d4"),
  3218 => (x"78",x"78",x"c0",x"78"),
  3219 => (x"c8",x"78",x"78",x"78"),
  3220 => (x"c7",x"c4",x"1e",x"c0"),
  3221 => (x"fb",x"fc",x"49",x"da"),
  3222 => (x"d0",x"ff",x"87",x"f7"),
  3223 => (x"c4",x"78",x"c4",x"48"),
  3224 => (x"d4",x"1e",x"da",x"c7"),
  3225 => (x"de",x"fd",x"49",x"66"),
  3226 => (x"1e",x"c1",x"87",x"ff"),
  3227 => (x"fd",x"49",x"66",x"d8"),
  3228 => (x"cc",x"87",x"cd",x"dc"),
  3229 => (x"48",x"66",x"dc",x"86"),
  3230 => (x"e0",x"c0",x"80",x"c1"),
  3231 => (x"ab",x"c1",x"58",x"a6"),
  3232 => (x"87",x"f3",x"c0",x"02"),
  3233 => (x"c1",x"49",x"66",x"cc"),
  3234 => (x"66",x"d0",x"81",x"d0"),
  3235 => (x"05",x"a8",x"69",x"48"),
  3236 => (x"a6",x"d0",x"87",x"dd"),
  3237 => (x"85",x"78",x"c1",x"48"),
  3238 => (x"c1",x"49",x"66",x"cc"),
  3239 => (x"ad",x"69",x"81",x"cc"),
  3240 => (x"c0",x"87",x"d4",x"05"),
  3241 => (x"48",x"66",x"d4",x"4d"),
  3242 => (x"a6",x"d8",x"80",x"c1"),
  3243 => (x"d0",x"87",x"c8",x"58"),
  3244 => (x"80",x"c1",x"48",x"66"),
  3245 => (x"c1",x"58",x"a6",x"d4"),
  3246 => (x"fd",x"05",x"8c",x"8b"),
  3247 => (x"66",x"d8",x"87",x"eb"),
  3248 => (x"dc",x"87",x"da",x"02"),
  3249 => (x"ff",x"c3",x"49",x"66"),
  3250 => (x"59",x"a6",x"d4",x"99"),
  3251 => (x"c8",x"49",x"66",x"dc"),
  3252 => (x"a6",x"d8",x"29",x"b7"),
  3253 => (x"49",x"66",x"dc",x"59"),
  3254 => (x"71",x"29",x"b7",x"d8"),
  3255 => (x"bf",x"97",x"6e",x"4d"),
  3256 => (x"99",x"f0",x"c3",x"49"),
  3257 => (x"1e",x"71",x"b1",x"75"),
  3258 => (x"c8",x"49",x"66",x"d8"),
  3259 => (x"1e",x"71",x"29",x"b7"),
  3260 => (x"dc",x"1e",x"66",x"dc"),
  3261 => (x"66",x"d4",x"1e",x"66"),
  3262 => (x"1e",x"49",x"bf",x"97"),
  3263 => (x"f3",x"ea",x"49",x"c0"),
  3264 => (x"73",x"86",x"d4",x"87"),
  3265 => (x"87",x"c7",x"02",x"9b"),
  3266 => (x"cf",x"e2",x"49",x"d0"),
  3267 => (x"c2",x"87",x"c6",x"87"),
  3268 => (x"c7",x"e2",x"49",x"d0"),
  3269 => (x"05",x"9b",x"73",x"87"),
  3270 => (x"e0",x"87",x"e1",x"fb"),
  3271 => (x"87",x"d5",x"e3",x"8e"),
  3272 => (x"5c",x"5b",x"5e",x"0e"),
  3273 => (x"86",x"e4",x"0e",x"5d"),
  3274 => (x"a6",x"cc",x"4a",x"71"),
  3275 => (x"78",x"ff",x"c0",x"48"),
  3276 => (x"ff",x"c1",x"80",x"c4"),
  3277 => (x"c3",x"80",x"c4",x"78"),
  3278 => (x"80",x"c4",x"78",x"ff"),
  3279 => (x"a2",x"c8",x"78",x"c0"),
  3280 => (x"c9",x"49",x"69",x"49"),
  3281 => (x"9d",x"4d",x"71",x"29"),
  3282 => (x"87",x"ee",x"c2",x"02"),
  3283 => (x"a6",x"cc",x"4c",x"c0"),
  3284 => (x"c2",x"02",x"6b",x"4b"),
  3285 => (x"49",x"74",x"87",x"ca"),
  3286 => (x"a1",x"73",x"91",x"c4"),
  3287 => (x"c8",x"7e",x"69",x"49"),
  3288 => (x"78",x"c4",x"48",x"a6"),
  3289 => (x"6e",x"49",x"66",x"c8"),
  3290 => (x"72",x"1e",x"71",x"91"),
  3291 => (x"4a",x"09",x"75",x"1e"),
  3292 => (x"87",x"c5",x"f6",x"fc"),
  3293 => (x"49",x"26",x"4a",x"26"),
  3294 => (x"c4",x"58",x"a6",x"c8"),
  3295 => (x"b7",x"c0",x"c0",x"c0"),
  3296 => (x"87",x"cb",x"01",x"ad"),
  3297 => (x"a8",x"b7",x"ff",x"cf"),
  3298 => (x"87",x"fd",x"c0",x"06"),
  3299 => (x"c4",x"87",x"eb",x"c0"),
  3300 => (x"ff",x"c3",x"48",x"66"),
  3301 => (x"04",x"a8",x"b7",x"ff"),
  3302 => (x"c4",x"87",x"ee",x"c0"),
  3303 => (x"ff",x"c7",x"48",x"66"),
  3304 => (x"03",x"a8",x"b7",x"ff"),
  3305 => (x"66",x"c8",x"87",x"c9"),
  3306 => (x"a8",x"b7",x"c5",x"48"),
  3307 => (x"c4",x"87",x"da",x"03"),
  3308 => (x"ff",x"cf",x"48",x"66"),
  3309 => (x"06",x"a8",x"b7",x"ff"),
  3310 => (x"66",x"c8",x"87",x"cf"),
  3311 => (x"cc",x"80",x"c1",x"48"),
  3312 => (x"b7",x"d0",x"58",x"a6"),
  3313 => (x"db",x"fe",x"06",x"a8"),
  3314 => (x"48",x"66",x"c8",x"87"),
  3315 => (x"06",x"a8",x"b7",x"d0"),
  3316 => (x"84",x"c1",x"87",x"ce"),
  3317 => (x"91",x"c4",x"49",x"74"),
  3318 => (x"69",x"49",x"a1",x"73"),
  3319 => (x"87",x"f6",x"fd",x"05"),
  3320 => (x"49",x"a2",x"c8",x"c1"),
  3321 => (x"c1",x"79",x"66",x"c4"),
  3322 => (x"c8",x"49",x"a2",x"cc"),
  3323 => (x"d0",x"c1",x"79",x"66"),
  3324 => (x"79",x"6e",x"49",x"a2"),
  3325 => (x"49",x"a2",x"d4",x"c1"),
  3326 => (x"8e",x"e4",x"79",x"c1"),
  3327 => (x"87",x"f5",x"df",x"ff"),
  3328 => (x"c4",x"49",x"c0",x"1e"),
  3329 => (x"02",x"bf",x"eb",x"dc"),
  3330 => (x"49",x"c1",x"87",x"c2"),
  3331 => (x"bf",x"c7",x"de",x"c4"),
  3332 => (x"c2",x"87",x"c2",x"02"),
  3333 => (x"48",x"d0",x"ff",x"b1"),
  3334 => (x"ff",x"78",x"c5",x"c8"),
  3335 => (x"fa",x"c3",x"48",x"d4"),
  3336 => (x"ff",x"78",x"71",x"78"),
  3337 => (x"78",x"c4",x"48",x"d0"),
  3338 => (x"73",x"1e",x"4f",x"26"),
  3339 => (x"1e",x"4a",x"71",x"1e"),
  3340 => (x"c1",x"49",x"66",x"cc"),
  3341 => (x"dc",x"c4",x"91",x"dc"),
  3342 => (x"83",x"71",x"4b",x"e3"),
  3343 => (x"d0",x"fd",x"49",x"73"),
  3344 => (x"86",x"c4",x"87",x"f1"),
  3345 => (x"c5",x"02",x"98",x"70"),
  3346 => (x"fb",x"49",x"73",x"87"),
  3347 => (x"ef",x"fe",x"87",x"d2"),
  3348 => (x"e4",x"de",x"ff",x"87"),
  3349 => (x"5b",x"5e",x"0e",x"87"),
  3350 => (x"f4",x"0e",x"5d",x"5c"),
  3351 => (x"d3",x"dd",x"ff",x"86"),
  3352 => (x"c4",x"49",x"70",x"87"),
  3353 => (x"d2",x"c5",x"02",x"99"),
  3354 => (x"48",x"d0",x"ff",x"87"),
  3355 => (x"ff",x"78",x"c5",x"c8"),
  3356 => (x"c0",x"c2",x"48",x"d4"),
  3357 => (x"78",x"78",x"c0",x"78"),
  3358 => (x"4d",x"78",x"78",x"78"),
  3359 => (x"c0",x"48",x"d4",x"ff"),
  3360 => (x"a5",x"4a",x"76",x"78"),
  3361 => (x"bf",x"d4",x"ff",x"49"),
  3362 => (x"d4",x"ff",x"79",x"97"),
  3363 => (x"68",x"78",x"c0",x"48"),
  3364 => (x"c8",x"85",x"c1",x"51"),
  3365 => (x"e3",x"04",x"ad",x"b7"),
  3366 => (x"48",x"d0",x"ff",x"87"),
  3367 => (x"97",x"c6",x"78",x"c4"),
  3368 => (x"a6",x"cc",x"48",x"66"),
  3369 => (x"d0",x"4c",x"70",x"58"),
  3370 => (x"2c",x"b7",x"c4",x"9c"),
  3371 => (x"dc",x"c1",x"49",x"74"),
  3372 => (x"e3",x"dc",x"c4",x"91"),
  3373 => (x"69",x"81",x"c8",x"81"),
  3374 => (x"c2",x"87",x"ca",x"05"),
  3375 => (x"db",x"ff",x"49",x"d1"),
  3376 => (x"f6",x"c3",x"87",x"da"),
  3377 => (x"66",x"97",x"c7",x"87"),
  3378 => (x"f0",x"c3",x"49",x"4b"),
  3379 => (x"05",x"a9",x"d0",x"99"),
  3380 => (x"1e",x"74",x"87",x"cc"),
  3381 => (x"d2",x"e4",x"49",x"72"),
  3382 => (x"c3",x"86",x"c4",x"87"),
  3383 => (x"d0",x"c2",x"87",x"dd"),
  3384 => (x"87",x"c8",x"05",x"ab"),
  3385 => (x"e5",x"e4",x"49",x"72"),
  3386 => (x"87",x"cf",x"c3",x"87"),
  3387 => (x"05",x"ab",x"ec",x"c3"),
  3388 => (x"1e",x"c0",x"87",x"ce"),
  3389 => (x"49",x"72",x"1e",x"74"),
  3390 => (x"c8",x"87",x"cf",x"e5"),
  3391 => (x"87",x"fb",x"c2",x"86"),
  3392 => (x"05",x"ab",x"d1",x"c2"),
  3393 => (x"1e",x"74",x"87",x"cc"),
  3394 => (x"ea",x"e6",x"49",x"72"),
  3395 => (x"c2",x"86",x"c4",x"87"),
  3396 => (x"c6",x"c3",x"87",x"e9"),
  3397 => (x"87",x"cc",x"05",x"ab"),
  3398 => (x"49",x"72",x"1e",x"74"),
  3399 => (x"c4",x"87",x"cd",x"e7"),
  3400 => (x"87",x"d7",x"c2",x"86"),
  3401 => (x"05",x"ab",x"e0",x"c0"),
  3402 => (x"1e",x"c0",x"87",x"ce"),
  3403 => (x"49",x"72",x"1e",x"74"),
  3404 => (x"c8",x"87",x"e5",x"e9"),
  3405 => (x"87",x"c3",x"c2",x"86"),
  3406 => (x"05",x"ab",x"c4",x"c3"),
  3407 => (x"1e",x"c1",x"87",x"ce"),
  3408 => (x"49",x"72",x"1e",x"74"),
  3409 => (x"c8",x"87",x"d1",x"e9"),
  3410 => (x"87",x"ef",x"c1",x"86"),
  3411 => (x"05",x"ab",x"f0",x"c0"),
  3412 => (x"1e",x"c0",x"87",x"ce"),
  3413 => (x"49",x"72",x"1e",x"74"),
  3414 => (x"c8",x"87",x"d0",x"f0"),
  3415 => (x"87",x"db",x"c1",x"86"),
  3416 => (x"05",x"ab",x"c5",x"c3"),
  3417 => (x"1e",x"c1",x"87",x"ce"),
  3418 => (x"49",x"72",x"1e",x"74"),
  3419 => (x"c8",x"87",x"fc",x"ef"),
  3420 => (x"87",x"c7",x"c1",x"86"),
  3421 => (x"cc",x"05",x"ab",x"c8"),
  3422 => (x"72",x"1e",x"74",x"87"),
  3423 => (x"87",x"c7",x"e7",x"49"),
  3424 => (x"f6",x"c0",x"86",x"c4"),
  3425 => (x"05",x"9b",x"73",x"87"),
  3426 => (x"1e",x"74",x"87",x"cc"),
  3427 => (x"fb",x"e5",x"49",x"72"),
  3428 => (x"c0",x"86",x"c4",x"87"),
  3429 => (x"66",x"c8",x"87",x"e5"),
  3430 => (x"66",x"97",x"c9",x"1e"),
  3431 => (x"97",x"cc",x"1e",x"49"),
  3432 => (x"cf",x"1e",x"49",x"66"),
  3433 => (x"1e",x"49",x"66",x"97"),
  3434 => (x"49",x"66",x"97",x"d2"),
  3435 => (x"e0",x"49",x"c4",x"1e"),
  3436 => (x"86",x"d4",x"87",x"c2"),
  3437 => (x"ff",x"49",x"d1",x"c2"),
  3438 => (x"f4",x"87",x"e1",x"d7"),
  3439 => (x"f4",x"d8",x"ff",x"8e"),
  3440 => (x"d8",x"c3",x"1e",x"87"),
  3441 => (x"c1",x"49",x"bf",x"cf"),
  3442 => (x"d3",x"d8",x"c3",x"b9"),
  3443 => (x"48",x"d4",x"ff",x"59"),
  3444 => (x"ff",x"78",x"ff",x"c3"),
  3445 => (x"e1",x"c0",x"48",x"d0"),
  3446 => (x"48",x"d4",x"ff",x"78"),
  3447 => (x"31",x"c4",x"78",x"c1"),
  3448 => (x"d0",x"ff",x"78",x"71"),
  3449 => (x"78",x"e0",x"c0",x"48"),
  3450 => (x"c3",x"1e",x"4f",x"26"),
  3451 => (x"c4",x"1e",x"c3",x"d8"),
  3452 => (x"fd",x"49",x"d0",x"d4"),
  3453 => (x"c4",x"87",x"fc",x"c9"),
  3454 => (x"02",x"98",x"70",x"86"),
  3455 => (x"c0",x"ff",x"87",x"c3"),
  3456 => (x"31",x"4f",x"26",x"87"),
  3457 => (x"5a",x"48",x"4b",x"35"),
  3458 => (x"43",x"20",x"20",x"20"),
  3459 => (x"00",x"00",x"47",x"46"),
  3460 => (x"1e",x"00",x"00",x"00"),
  3461 => (x"87",x"de",x"c1",x"ff"),
  3462 => (x"87",x"c6",x"d5",x"fe"),
  3463 => (x"c2",x"49",x"66",x"c4"),
  3464 => (x"cd",x"02",x"99",x"c0"),
  3465 => (x"1e",x"e0",x"c3",x"87"),
  3466 => (x"49",x"fe",x"d8",x"c4"),
  3467 => (x"87",x"d7",x"d8",x"fe"),
  3468 => (x"66",x"c4",x"86",x"c4"),
  3469 => (x"99",x"c0",x"c4",x"49"),
  3470 => (x"c3",x"87",x"cd",x"02"),
  3471 => (x"d8",x"c4",x"1e",x"f0"),
  3472 => (x"d8",x"fe",x"49",x"fe"),
  3473 => (x"86",x"c4",x"87",x"c1"),
  3474 => (x"c1",x"49",x"66",x"c4"),
  3475 => (x"1e",x"71",x"99",x"ff"),
  3476 => (x"49",x"fe",x"d8",x"c4"),
  3477 => (x"87",x"ef",x"d7",x"fe"),
  3478 => (x"87",x"fe",x"d3",x"fe"),
  3479 => (x"0e",x"4f",x"26",x"26"),
  3480 => (x"5d",x"5c",x"5b",x"5e"),
  3481 => (x"86",x"d8",x"ff",x"0e"),
  3482 => (x"df",x"c4",x"7e",x"c0"),
  3483 => (x"c2",x"49",x"bf",x"df"),
  3484 => (x"72",x"1e",x"71",x"81"),
  3485 => (x"fc",x"4a",x"c6",x"1e"),
  3486 => (x"71",x"87",x"fe",x"e9"),
  3487 => (x"26",x"4a",x"26",x"48"),
  3488 => (x"58",x"a6",x"c8",x"49"),
  3489 => (x"bf",x"df",x"df",x"c4"),
  3490 => (x"71",x"81",x"c4",x"49"),
  3491 => (x"c6",x"1e",x"72",x"1e"),
  3492 => (x"e4",x"e9",x"fc",x"4a"),
  3493 => (x"26",x"48",x"71",x"87"),
  3494 => (x"cc",x"49",x"26",x"4a"),
  3495 => (x"e4",x"c3",x"58",x"a6"),
  3496 => (x"ff",x"49",x"bf",x"f2"),
  3497 => (x"70",x"87",x"d2",x"cc"),
  3498 => (x"fa",x"c9",x"02",x"98"),
  3499 => (x"49",x"e0",x"c0",x"87"),
  3500 => (x"87",x"f9",x"cb",x"ff"),
  3501 => (x"e4",x"c3",x"49",x"70"),
  3502 => (x"4c",x"c0",x"59",x"f6"),
  3503 => (x"91",x"c4",x"49",x"74"),
  3504 => (x"69",x"81",x"d0",x"fe"),
  3505 => (x"c4",x"49",x"74",x"4a"),
  3506 => (x"81",x"bf",x"df",x"df"),
  3507 => (x"df",x"c4",x"91",x"c4"),
  3508 => (x"79",x"72",x"81",x"eb"),
  3509 => (x"87",x"d2",x"02",x"9a"),
  3510 => (x"89",x"c1",x"49",x"72"),
  3511 => (x"48",x"6e",x"9a",x"71"),
  3512 => (x"7e",x"70",x"80",x"c1"),
  3513 => (x"ff",x"05",x"9a",x"72"),
  3514 => (x"84",x"c1",x"87",x"ee"),
  3515 => (x"04",x"ac",x"b7",x"c2"),
  3516 => (x"6e",x"87",x"c9",x"ff"),
  3517 => (x"b7",x"fc",x"c0",x"48"),
  3518 => (x"ea",x"c8",x"04",x"a8"),
  3519 => (x"74",x"4c",x"c0",x"87"),
  3520 => (x"82",x"66",x"c4",x"4a"),
  3521 => (x"df",x"c4",x"92",x"c4"),
  3522 => (x"49",x"74",x"82",x"eb"),
  3523 => (x"c4",x"81",x"66",x"c8"),
  3524 => (x"eb",x"df",x"c4",x"91"),
  3525 => (x"69",x"4a",x"6a",x"81"),
  3526 => (x"74",x"b9",x"72",x"49"),
  3527 => (x"df",x"df",x"c4",x"4b"),
  3528 => (x"93",x"c4",x"83",x"bf"),
  3529 => (x"83",x"eb",x"df",x"c4"),
  3530 => (x"48",x"72",x"ba",x"6b"),
  3531 => (x"a6",x"d4",x"98",x"71"),
  3532 => (x"c4",x"49",x"74",x"58"),
  3533 => (x"81",x"bf",x"df",x"df"),
  3534 => (x"df",x"c4",x"91",x"c4"),
  3535 => (x"7e",x"69",x"81",x"eb"),
  3536 => (x"c0",x"48",x"a6",x"d4"),
  3537 => (x"5c",x"a6",x"d0",x"78"),
  3538 => (x"d0",x"4c",x"ff",x"c3"),
  3539 => (x"29",x"df",x"49",x"66"),
  3540 => (x"87",x"e2",x"c6",x"02"),
  3541 => (x"c0",x"4a",x"66",x"cc"),
  3542 => (x"66",x"d4",x"92",x"e0"),
  3543 => (x"48",x"ff",x"c0",x"82"),
  3544 => (x"4a",x"70",x"88",x"72"),
  3545 => (x"c0",x"48",x"a6",x"d8"),
  3546 => (x"c0",x"80",x"c4",x"78"),
  3547 => (x"df",x"49",x"6e",x"78"),
  3548 => (x"a6",x"e4",x"c0",x"29"),
  3549 => (x"db",x"df",x"c4",x"59"),
  3550 => (x"72",x"78",x"c1",x"48"),
  3551 => (x"b7",x"31",x"c3",x"49"),
  3552 => (x"c0",x"b1",x"72",x"2a"),
  3553 => (x"91",x"c4",x"99",x"ff"),
  3554 => (x"4d",x"c8",x"c0",x"c4"),
  3555 => (x"4b",x"6d",x"85",x"71"),
  3556 => (x"c0",x"c0",x"c4",x"49"),
  3557 => (x"87",x"d7",x"02",x"99"),
  3558 => (x"02",x"66",x"e0",x"c0"),
  3559 => (x"c8",x"87",x"c7",x"c0"),
  3560 => (x"c5",x"78",x"c0",x"80"),
  3561 => (x"df",x"c4",x"87",x"d0"),
  3562 => (x"78",x"c1",x"48",x"e3"),
  3563 => (x"c0",x"87",x"c7",x"c5"),
  3564 => (x"d8",x"02",x"66",x"e0"),
  3565 => (x"c2",x"49",x"73",x"87"),
  3566 => (x"02",x"99",x"c0",x"c0"),
  3567 => (x"d0",x"87",x"c3",x"c0"),
  3568 => (x"48",x"6d",x"2b",x"b7"),
  3569 => (x"98",x"ff",x"ff",x"fd"),
  3570 => (x"fa",x"c0",x"7d",x"70"),
  3571 => (x"e3",x"df",x"c4",x"87"),
  3572 => (x"f2",x"c0",x"02",x"bf"),
  3573 => (x"d0",x"48",x"73",x"87"),
  3574 => (x"e8",x"c0",x"28",x"b7"),
  3575 => (x"98",x"70",x"58",x"a6"),
  3576 => (x"87",x"e3",x"c0",x"02"),
  3577 => (x"bf",x"e7",x"df",x"c4"),
  3578 => (x"c0",x"e0",x"c0",x"49"),
  3579 => (x"ca",x"c0",x"02",x"99"),
  3580 => (x"c0",x"49",x"70",x"87"),
  3581 => (x"02",x"99",x"c0",x"e0"),
  3582 => (x"6d",x"87",x"cc",x"c0"),
  3583 => (x"c0",x"c0",x"c2",x"48"),
  3584 => (x"c0",x"7d",x"70",x"b0"),
  3585 => (x"73",x"4b",x"66",x"e4"),
  3586 => (x"c0",x"c0",x"c8",x"49"),
  3587 => (x"c5",x"c2",x"02",x"99"),
  3588 => (x"e7",x"df",x"c4",x"87"),
  3589 => (x"c0",x"cc",x"4a",x"bf"),
  3590 => (x"cf",x"c0",x"02",x"9a"),
  3591 => (x"8a",x"c0",x"c4",x"87"),
  3592 => (x"87",x"d7",x"c0",x"02"),
  3593 => (x"f8",x"c0",x"02",x"8a"),
  3594 => (x"87",x"dc",x"c1",x"87"),
  3595 => (x"99",x"74",x"49",x"73"),
  3596 => (x"ff",x"c3",x"91",x"c2"),
  3597 => (x"4b",x"11",x"81",x"fc"),
  3598 => (x"73",x"87",x"db",x"c1"),
  3599 => (x"c2",x"99",x"74",x"49"),
  3600 => (x"fc",x"ff",x"c3",x"91"),
  3601 => (x"11",x"81",x"c1",x"81"),
  3602 => (x"66",x"e0",x"c0",x"4b"),
  3603 => (x"87",x"c8",x"c0",x"02"),
  3604 => (x"d2",x"48",x"a6",x"dc"),
  3605 => (x"87",x"fe",x"c0",x"78"),
  3606 => (x"c4",x"48",x"a6",x"d8"),
  3607 => (x"f5",x"c0",x"78",x"d2"),
  3608 => (x"74",x"49",x"73",x"87"),
  3609 => (x"c3",x"91",x"c2",x"99"),
  3610 => (x"c1",x"81",x"fc",x"ff"),
  3611 => (x"c0",x"4b",x"11",x"81"),
  3612 => (x"c0",x"02",x"66",x"e0"),
  3613 => (x"a6",x"dc",x"87",x"c9"),
  3614 => (x"78",x"d9",x"c1",x"48"),
  3615 => (x"d8",x"87",x"d7",x"c0"),
  3616 => (x"d9",x"c5",x"48",x"a6"),
  3617 => (x"87",x"ce",x"c0",x"78"),
  3618 => (x"99",x"74",x"49",x"73"),
  3619 => (x"ff",x"c3",x"91",x"c2"),
  3620 => (x"81",x"c1",x"81",x"fc"),
  3621 => (x"e0",x"c0",x"4b",x"11"),
  3622 => (x"db",x"c0",x"02",x"66"),
  3623 => (x"ff",x"49",x"73",x"87"),
  3624 => (x"c0",x"fc",x"c7",x"b9"),
  3625 => (x"c4",x"48",x"71",x"99"),
  3626 => (x"98",x"bf",x"e7",x"df"),
  3627 => (x"58",x"eb",x"df",x"c4"),
  3628 => (x"c0",x"c4",x"9b",x"74"),
  3629 => (x"87",x"d3",x"c0",x"b3"),
  3630 => (x"fc",x"c7",x"49",x"73"),
  3631 => (x"48",x"71",x"99",x"c0"),
  3632 => (x"bf",x"e7",x"df",x"c4"),
  3633 => (x"eb",x"df",x"c4",x"b0"),
  3634 => (x"d8",x"9b",x"74",x"58"),
  3635 => (x"ca",x"c0",x"02",x"66"),
  3636 => (x"df",x"c4",x"1e",x"87"),
  3637 => (x"fa",x"f4",x"49",x"db"),
  3638 => (x"73",x"86",x"c4",x"87"),
  3639 => (x"db",x"df",x"c4",x"1e"),
  3640 => (x"87",x"ef",x"f4",x"49"),
  3641 => (x"66",x"dc",x"86",x"c4"),
  3642 => (x"87",x"ca",x"c0",x"02"),
  3643 => (x"db",x"df",x"c4",x"1e"),
  3644 => (x"87",x"df",x"f4",x"49"),
  3645 => (x"66",x"d0",x"86",x"c4"),
  3646 => (x"d4",x"30",x"c1",x"48"),
  3647 => (x"48",x"6e",x"58",x"a6"),
  3648 => (x"7e",x"70",x"30",x"c1"),
  3649 => (x"c1",x"48",x"66",x"d4"),
  3650 => (x"58",x"a6",x"d8",x"80"),
  3651 => (x"a8",x"b7",x"e0",x"c0"),
  3652 => (x"87",x"f7",x"f8",x"04"),
  3653 => (x"c1",x"4c",x"66",x"cc"),
  3654 => (x"ac",x"b7",x"c2",x"84"),
  3655 => (x"87",x"df",x"f7",x"04"),
  3656 => (x"48",x"df",x"df",x"c4"),
  3657 => (x"ff",x"78",x"66",x"c4"),
  3658 => (x"4d",x"26",x"8e",x"d8"),
  3659 => (x"4b",x"26",x"4c",x"26"),
  3660 => (x"00",x"00",x"4f",x"26"),
  3661 => (x"c0",x"1e",x"00",x"00"),
  3662 => (x"c4",x"49",x"72",x"4a"),
  3663 => (x"eb",x"df",x"c4",x"91"),
  3664 => (x"c1",x"79",x"ff",x"81"),
  3665 => (x"aa",x"b7",x"c6",x"82"),
  3666 => (x"c4",x"87",x"ee",x"04"),
  3667 => (x"c0",x"48",x"df",x"df"),
  3668 => (x"26",x"78",x"40",x"40"),
  3669 => (x"71",x"1e",x"1e",x"4f"),
  3670 => (x"c7",x"e0",x"c4",x"4a"),
  3671 => (x"c1",x"48",x"7e",x"bf"),
  3672 => (x"cb",x"e0",x"c4",x"80"),
  3673 => (x"81",x"c4",x"49",x"58"),
  3674 => (x"51",x"72",x"81",x"6e"),
  3675 => (x"e0",x"c4",x"98",x"cf"),
  3676 => (x"dc",x"48",x"58",x"cb"),
  3677 => (x"c8",x"40",x"c6",x"80"),
  3678 => (x"66",x"cc",x"78",x"66"),
  3679 => (x"ec",x"c0",x"ff",x"49"),
  3680 => (x"c4",x"49",x"70",x"87"),
  3681 => (x"26",x"59",x"e3",x"e0"),
  3682 => (x"73",x"1e",x"4f",x"26"),
  3683 => (x"49",x"4a",x"71",x"1e"),
  3684 => (x"c0",x"02",x"99",x"c1"),
  3685 => (x"66",x"c8",x"87",x"eb"),
  3686 => (x"02",x"99",x"c1",x"49"),
  3687 => (x"c0",x"c3",x"87",x"c5"),
  3688 => (x"c3",x"87",x"c3",x"4b"),
  3689 => (x"c8",x"c3",x"4b",x"d0"),
  3690 => (x"73",x"1e",x"c4",x"1e"),
  3691 => (x"fe",x"b1",x"c7",x"49"),
  3692 => (x"c8",x"c3",x"87",x"e3"),
  3693 => (x"dc",x"1e",x"c4",x"1e"),
  3694 => (x"b1",x"73",x"49",x"66"),
  3695 => (x"d0",x"87",x"d6",x"fe"),
  3696 => (x"87",x"ea",x"fd",x"86"),
  3697 => (x"5c",x"5b",x"5e",x"0e"),
  3698 => (x"86",x"f8",x"0e",x"5d"),
  3699 => (x"bf",x"df",x"e0",x"c4"),
  3700 => (x"e4",x"ff",x"fe",x"49"),
  3701 => (x"7e",x"49",x"70",x"87"),
  3702 => (x"db",x"fe",x"49",x"c4"),
  3703 => (x"d4",x"ff",x"87",x"ea"),
  3704 => (x"78",x"ff",x"c3",x"48"),
  3705 => (x"ff",x"c3",x"49",x"68"),
  3706 => (x"48",x"a6",x"c4",x"78"),
  3707 => (x"78",x"bf",x"d4",x"ff"),
  3708 => (x"c0",x"48",x"d0",x"ff"),
  3709 => (x"e1",x"c2",x"78",x"e0"),
  3710 => (x"f1",x"c2",x"05",x"a9"),
  3711 => (x"4a",x"66",x"c4",x"87"),
  3712 => (x"02",x"8a",x"e0",x"c0"),
  3713 => (x"d0",x"87",x"c3",x"c2"),
  3714 => (x"d3",x"c2",x"02",x"8a"),
  3715 => (x"02",x"8a",x"c1",x"87"),
  3716 => (x"8a",x"87",x"cd",x"c2"),
  3717 => (x"87",x"c8",x"c2",x"02"),
  3718 => (x"c3",x"c2",x"02",x"8a"),
  3719 => (x"02",x"8a",x"cc",x"87"),
  3720 => (x"c2",x"87",x"f5",x"c1"),
  3721 => (x"c0",x"02",x"8a",x"fe"),
  3722 => (x"8a",x"c1",x"87",x"fd"),
  3723 => (x"8a",x"87",x"d5",x"02"),
  3724 => (x"87",x"fa",x"c1",x"05"),
  3725 => (x"c1",x"1e",x"c8",x"c3"),
  3726 => (x"49",x"ff",x"c3",x"1e"),
  3727 => (x"c8",x"87",x"d6",x"fc"),
  3728 => (x"87",x"ea",x"c1",x"86"),
  3729 => (x"bf",x"e3",x"e0",x"c4"),
  3730 => (x"05",x"a8",x"c1",x"48"),
  3731 => (x"c8",x"c3",x"87",x"d0"),
  3732 => (x"c3",x"1e",x"c2",x"1e"),
  3733 => (x"fc",x"fb",x"49",x"fe"),
  3734 => (x"c1",x"86",x"c8",x"87"),
  3735 => (x"e0",x"c4",x"87",x"d0"),
  3736 => (x"78",x"c0",x"48",x"e3"),
  3737 => (x"c4",x"87",x"c7",x"c1"),
  3738 => (x"48",x"bf",x"e3",x"e0"),
  3739 => (x"d0",x"05",x"a8",x"c2"),
  3740 => (x"1e",x"c8",x"c3",x"87"),
  3741 => (x"fd",x"c3",x"1e",x"c3"),
  3742 => (x"87",x"d9",x"fb",x"49"),
  3743 => (x"ed",x"c0",x"86",x"c8"),
  3744 => (x"e3",x"e0",x"c4",x"87"),
  3745 => (x"c0",x"78",x"c0",x"48"),
  3746 => (x"1e",x"c0",x"87",x"e4"),
  3747 => (x"c1",x"c2",x"1e",x"c3"),
  3748 => (x"87",x"c1",x"fb",x"49"),
  3749 => (x"87",x"d6",x"86",x"c8"),
  3750 => (x"48",x"e3",x"e0",x"c4"),
  3751 => (x"87",x"ce",x"78",x"c3"),
  3752 => (x"c3",x"48",x"66",x"c4"),
  3753 => (x"df",x"e0",x"c4",x"98"),
  3754 => (x"80",x"c8",x"48",x"58"),
  3755 => (x"e0",x"c4",x"78",x"c3"),
  3756 => (x"c2",x"4b",x"bf",x"e3"),
  3757 => (x"e4",x"c0",x"02",x"8b"),
  3758 => (x"02",x"8b",x"c1",x"87"),
  3759 => (x"8b",x"87",x"f3",x"c0"),
  3760 => (x"8b",x"87",x"cc",x"02"),
  3761 => (x"8b",x"87",x"c8",x"02"),
  3762 => (x"87",x"ea",x"c3",x"02"),
  3763 => (x"6e",x"87",x"e5",x"c4"),
  3764 => (x"87",x"e0",x"c4",x"02"),
  3765 => (x"48",x"e3",x"e0",x"c4"),
  3766 => (x"d7",x"c4",x"78",x"c3"),
  3767 => (x"c4",x"02",x"6e",x"87"),
  3768 => (x"c8",x"c3",x"87",x"d2"),
  3769 => (x"c3",x"1e",x"c1",x"1e"),
  3770 => (x"e8",x"f9",x"49",x"ff"),
  3771 => (x"c4",x"86",x"c8",x"87"),
  3772 => (x"e0",x"c4",x"87",x"c2"),
  3773 => (x"c2",x"49",x"bf",x"db"),
  3774 => (x"f3",x"c1",x"02",x"99"),
  3775 => (x"eb",x"e0",x"c4",x"87"),
  3776 => (x"c8",x"c0",x"05",x"bf"),
  3777 => (x"ef",x"e0",x"c4",x"87"),
  3778 => (x"e3",x"c1",x"02",x"bf"),
  3779 => (x"eb",x"e0",x"c4",x"87"),
  3780 => (x"ff",x"4c",x"4d",x"bf"),
  3781 => (x"03",x"ad",x"b7",x"c0"),
  3782 => (x"4c",x"87",x"c1",x"c0"),
  3783 => (x"ac",x"b7",x"ff",x"c0"),
  3784 => (x"87",x"c1",x"c0",x"06"),
  3785 => (x"74",x"48",x"75",x"4c"),
  3786 => (x"ef",x"e0",x"c4",x"88"),
  3787 => (x"1e",x"c8",x"c3",x"58"),
  3788 => (x"49",x"74",x"1e",x"c4"),
  3789 => (x"f8",x"99",x"ff",x"c1"),
  3790 => (x"86",x"c8",x"87",x"db"),
  3791 => (x"bf",x"ef",x"e0",x"c4"),
  3792 => (x"8c",x"0c",x"c0",x"4c"),
  3793 => (x"ac",x"b7",x"c0",x"ff"),
  3794 => (x"87",x"c1",x"c0",x"03"),
  3795 => (x"b7",x"ff",x"c0",x"4c"),
  3796 => (x"c1",x"c0",x"06",x"ac"),
  3797 => (x"e0",x"c4",x"4c",x"87"),
  3798 => (x"74",x"48",x"bf",x"ef"),
  3799 => (x"f3",x"e0",x"c4",x"80"),
  3800 => (x"1e",x"c8",x"c3",x"58"),
  3801 => (x"49",x"74",x"1e",x"c5"),
  3802 => (x"f7",x"99",x"ff",x"c1"),
  3803 => (x"86",x"c8",x"87",x"e7"),
  3804 => (x"bf",x"db",x"e0",x"c4"),
  3805 => (x"02",x"99",x"c1",x"49"),
  3806 => (x"c4",x"87",x"fb",x"c0"),
  3807 => (x"4c",x"bf",x"f3",x"e0"),
  3808 => (x"bf",x"d0",x"f0",x"c3"),
  3809 => (x"c0",x"bb",x"74",x"4b"),
  3810 => (x"73",x"1e",x"74",x"1e"),
  3811 => (x"87",x"fa",x"f7",x"49"),
  3812 => (x"b7",x"2b",x"b7",x"c1"),
  3813 => (x"74",x"1e",x"c2",x"2c"),
  3814 => (x"f7",x"49",x"73",x"1e"),
  3815 => (x"b7",x"c1",x"87",x"ec"),
  3816 => (x"1e",x"2c",x"b7",x"2b"),
  3817 => (x"49",x"73",x"1e",x"74"),
  3818 => (x"d8",x"87",x"df",x"f7"),
  3819 => (x"d0",x"f0",x"c3",x"86"),
  3820 => (x"f3",x"e0",x"c4",x"48"),
  3821 => (x"e0",x"c4",x"78",x"bf"),
  3822 => (x"c4",x"48",x"bf",x"c7"),
  3823 => (x"a8",x"bf",x"c3",x"e0"),
  3824 => (x"87",x"f0",x"c0",x"02"),
  3825 => (x"80",x"c1",x"48",x"7e"),
  3826 => (x"58",x"c7",x"e0",x"c4"),
  3827 => (x"6e",x"83",x"c8",x"4b"),
  3828 => (x"4b",x"6b",x"97",x"83"),
  3829 => (x"e0",x"c4",x"98",x"cf"),
  3830 => (x"49",x"c5",x"58",x"c7"),
  3831 => (x"87",x"e8",x"d3",x"fe"),
  3832 => (x"73",x"48",x"d4",x"ff"),
  3833 => (x"48",x"d0",x"ff",x"78"),
  3834 => (x"c4",x"78",x"e0",x"c0"),
  3835 => (x"c4",x"48",x"e3",x"e0"),
  3836 => (x"78",x"bf",x"e7",x"e0"),
  3837 => (x"bf",x"c7",x"e0",x"c4"),
  3838 => (x"c3",x"e0",x"c4",x"48"),
  3839 => (x"c0",x"05",x"a8",x"bf"),
  3840 => (x"7e",x"c0",x"87",x"c5"),
  3841 => (x"c1",x"87",x"c2",x"c0"),
  3842 => (x"f8",x"48",x"6e",x"7e"),
  3843 => (x"87",x"da",x"f4",x"8e"),
  3844 => (x"00",x"00",x"00",x"00"),
  3845 => (x"5c",x"5b",x"5e",x"0e"),
  3846 => (x"4b",x"71",x"0e",x"5d"),
  3847 => (x"e0",x"c4",x"4c",x"c0"),
  3848 => (x"c4",x"05",x"bf",x"db"),
  3849 => (x"c2",x"4d",x"c1",x"87"),
  3850 => (x"75",x"4d",x"c0",x"87"),
  3851 => (x"05",x"99",x"c1",x"49"),
  3852 => (x"d0",x"87",x"e5",x"c1"),
  3853 => (x"87",x"c3",x"02",x"66"),
  3854 => (x"73",x"b3",x"c0",x"c2"),
  3855 => (x"ce",x"c9",x"fe",x"49"),
  3856 => (x"d4",x"4a",x"70",x"87"),
  3857 => (x"87",x"c6",x"05",x"66"),
  3858 => (x"c1",x"05",x"9a",x"72"),
  3859 => (x"fe",x"c3",x"87",x"ca"),
  3860 => (x"81",x"74",x"49",x"d3"),
  3861 => (x"02",x"9a",x"4a",x"11"),
  3862 => (x"73",x"87",x"fd",x"c0"),
  3863 => (x"f2",x"c0",x"05",x"aa"),
  3864 => (x"02",x"66",x"d4",x"87"),
  3865 => (x"d0",x"c3",x"87",x"c5"),
  3866 => (x"c3",x"87",x"c3",x"4d"),
  3867 => (x"c8",x"c3",x"4d",x"c0"),
  3868 => (x"74",x"1e",x"c4",x"1e"),
  3869 => (x"2a",x"b7",x"c4",x"4a"),
  3870 => (x"b1",x"75",x"49",x"72"),
  3871 => (x"c3",x"87",x"d6",x"f3"),
  3872 => (x"1e",x"c4",x"1e",x"c8"),
  3873 => (x"9a",x"cf",x"4a",x"74"),
  3874 => (x"b1",x"75",x"49",x"72"),
  3875 => (x"d0",x"87",x"c6",x"f3"),
  3876 => (x"c1",x"87",x"c5",x"86"),
  3877 => (x"87",x"f6",x"fe",x"84"),
  3878 => (x"1e",x"87",x"cf",x"f2"),
  3879 => (x"4b",x"71",x"1e",x"73"),
  3880 => (x"73",x"87",x"fc",x"e6"),
  3881 => (x"c1",x"c4",x"fe",x"49"),
  3882 => (x"87",x"c2",x"f2",x"87"),
  3883 => (x"fe",x"49",x"c1",x"1e"),
  3884 => (x"ff",x"87",x"d5",x"d0"),
  3885 => (x"d9",x"c4",x"48",x"d4"),
  3886 => (x"ff",x"78",x"bf",x"ea"),
  3887 => (x"e0",x"c0",x"48",x"d0"),
  3888 => (x"1e",x"4f",x"26",x"78"),
  3889 => (x"e0",x"c4",x"4a",x"c0"),
  3890 => (x"ca",x"02",x"bf",x"f7"),
  3891 => (x"e0",x"c4",x"49",x"87"),
  3892 => (x"a1",x"c1",x"48",x"f7"),
  3893 => (x"72",x"4a",x"11",x"78"),
  3894 => (x"87",x"c6",x"05",x"9a"),
  3895 => (x"48",x"f7",x"e0",x"c4"),
  3896 => (x"48",x"72",x"78",x"c0"),
  3897 => (x"c4",x"1e",x"4f",x"26"),
  3898 => (x"c4",x"48",x"f7",x"e0"),
  3899 => (x"78",x"bf",x"c8",x"c4"),
  3900 => (x"5e",x"0e",x"4f",x"26"),
  3901 => (x"0e",x"5d",x"5c",x"5b"),
  3902 => (x"c4",x"4b",x"71",x"1e"),
  3903 => (x"fd",x"49",x"d2",x"d9"),
  3904 => (x"70",x"87",x"f6",x"fb"),
  3905 => (x"d2",x"d9",x"c4",x"4d"),
  3906 => (x"ec",x"fb",x"fd",x"49"),
  3907 => (x"c4",x"7e",x"70",x"87"),
  3908 => (x"fd",x"49",x"d2",x"d9"),
  3909 => (x"70",x"87",x"e2",x"fb"),
  3910 => (x"05",x"ab",x"c4",x"4c"),
  3911 => (x"d9",x"c4",x"87",x"c8"),
  3912 => (x"fb",x"fd",x"49",x"d2"),
  3913 => (x"48",x"75",x"87",x"d3"),
  3914 => (x"e0",x"c4",x"98",x"c7"),
  3915 => (x"49",x"75",x"58",x"f7"),
  3916 => (x"02",x"99",x"e0",x"c0"),
  3917 => (x"49",x"74",x"87",x"c7"),
  3918 => (x"71",x"b1",x"c0",x"fc"),
  3919 => (x"d0",x"49",x"75",x"4c"),
  3920 => (x"87",x"c7",x"02",x"99"),
  3921 => (x"c0",x"fc",x"49",x"6e"),
  3922 => (x"c4",x"7e",x"71",x"b1"),
  3923 => (x"48",x"bf",x"eb",x"e0"),
  3924 => (x"e0",x"c4",x"80",x"6e"),
  3925 => (x"49",x"74",x"58",x"ef"),
  3926 => (x"c4",x"89",x"09",x"c0"),
  3927 => (x"48",x"bf",x"ef",x"e0"),
  3928 => (x"e0",x"c4",x"80",x"71"),
  3929 => (x"ef",x"26",x"58",x"f3"),
  3930 => (x"5e",x"0e",x"87",x"c0"),
  3931 => (x"0e",x"5d",x"5c",x"5b"),
  3932 => (x"ff",x"4d",x"d0",x"ff"),
  3933 => (x"c7",x"c4",x"4a",x"d4"),
  3934 => (x"7d",x"c5",x"4b",x"da"),
  3935 => (x"c3",x"7a",x"d5",x"c1"),
  3936 => (x"c3",x"7d",x"c4",x"7a"),
  3937 => (x"7d",x"c5",x"7a",x"ff"),
  3938 => (x"c3",x"7a",x"d7",x"c1"),
  3939 => (x"7d",x"c4",x"7a",x"ff"),
  3940 => (x"c1",x"7d",x"c5",x"c8"),
  3941 => (x"ff",x"c3",x"7a",x"d8"),
  3942 => (x"ff",x"c3",x"4c",x"7a"),
  3943 => (x"74",x"53",x"6a",x"7a"),
  3944 => (x"71",x"8c",x"c1",x"49"),
  3945 => (x"87",x"f2",x"05",x"99"),
  3946 => (x"7d",x"c5",x"7d",x"c4"),
  3947 => (x"c0",x"7a",x"d7",x"c1"),
  3948 => (x"ed",x"7d",x"c4",x"7a"),
  3949 => (x"5e",x"0e",x"87",x"f4"),
  3950 => (x"0e",x"5d",x"5c",x"5b"),
  3951 => (x"4d",x"c0",x"4b",x"71"),
  3952 => (x"c0",x"4c",x"66",x"d0"),
  3953 => (x"66",x"d0",x"8c",x"f0"),
  3954 => (x"87",x"ed",x"c0",x"02"),
  3955 => (x"02",x"8a",x"c3",x"4a"),
  3956 => (x"c0",x"87",x"e6",x"c0"),
  3957 => (x"c1",x"02",x"8a",x"ed"),
  3958 => (x"8a",x"c1",x"87",x"c4"),
  3959 => (x"87",x"fe",x"c0",x"02"),
  3960 => (x"db",x"c1",x"02",x"8a"),
  3961 => (x"c1",x"02",x"8a",x"87"),
  3962 => (x"8a",x"df",x"87",x"d6"),
  3963 => (x"87",x"e1",x"c1",x"02"),
  3964 => (x"c1",x"02",x"8a",x"c1"),
  3965 => (x"d5",x"c2",x"87",x"ee"),
  3966 => (x"02",x"9b",x"73",x"87"),
  3967 => (x"97",x"87",x"cf",x"c2"),
  3968 => (x"c9",x"c2",x"02",x"6b"),
  3969 => (x"ea",x"d9",x"c4",x"87"),
  3970 => (x"b0",x"c2",x"48",x"bf"),
  3971 => (x"58",x"ee",x"d9",x"c4"),
  3972 => (x"73",x"87",x"d9",x"fa"),
  3973 => (x"f3",x"c8",x"fd",x"49"),
  3974 => (x"c1",x"4d",x"70",x"87"),
  3975 => (x"1e",x"74",x"87",x"f0"),
  3976 => (x"f3",x"fe",x"49",x"c0"),
  3977 => (x"1e",x"74",x"87",x"f4"),
  3978 => (x"f3",x"fe",x"49",x"73"),
  3979 => (x"86",x"c8",x"87",x"ec"),
  3980 => (x"c8",x"c1",x"49",x"74"),
  3981 => (x"d3",x"da",x"c4",x"91"),
  3982 => (x"69",x"81",x"c8",x"81"),
  3983 => (x"87",x"ce",x"c1",x"4d"),
  3984 => (x"89",x"c2",x"49",x"74"),
  3985 => (x"49",x"73",x"1e",x"71"),
  3986 => (x"87",x"de",x"d7",x"ff"),
  3987 => (x"fd",x"c0",x"86",x"c4"),
  3988 => (x"cd",x"eb",x"c1",x"87"),
  3989 => (x"1e",x"50",x"c3",x"48"),
  3990 => (x"d9",x"fd",x"49",x"73"),
  3991 => (x"70",x"86",x"c4",x"87"),
  3992 => (x"87",x"ea",x"c0",x"4d"),
  3993 => (x"48",x"cd",x"eb",x"c1"),
  3994 => (x"1e",x"73",x"50",x"c3"),
  3995 => (x"49",x"d0",x"d4",x"c4"),
  3996 => (x"87",x"ff",x"e7",x"fc"),
  3997 => (x"98",x"70",x"86",x"c4"),
  3998 => (x"73",x"87",x"d3",x"02"),
  3999 => (x"87",x"ea",x"fb",x"49"),
  4000 => (x"1e",x"da",x"c7",x"c4"),
  4001 => (x"49",x"d0",x"d4",x"c4"),
  4002 => (x"87",x"dd",x"ee",x"fc"),
  4003 => (x"d9",x"c4",x"86",x"c4"),
  4004 => (x"fd",x"48",x"bf",x"ea"),
  4005 => (x"ee",x"d9",x"c4",x"98"),
  4006 => (x"87",x"d0",x"f8",x"58"),
  4007 => (x"c9",x"ea",x"48",x"75"),
  4008 => (x"1e",x"73",x"1e",x"87"),
  4009 => (x"d9",x"c4",x"4b",x"c0"),
  4010 => (x"78",x"c2",x"48",x"ea"),
  4011 => (x"48",x"c3",x"e0",x"c4"),
  4012 => (x"d4",x"78",x"40",x"c0"),
  4013 => (x"c8",x"78",x"c0",x"80"),
  4014 => (x"c1",x"78",x"c3",x"80"),
  4015 => (x"c0",x"48",x"cb",x"c1"),
  4016 => (x"87",x"e8",x"f7",x"50"),
  4017 => (x"48",x"cd",x"eb",x"c1"),
  4018 => (x"c3",x"1e",x"50",x"c3"),
  4019 => (x"fb",x"49",x"e4",x"fc"),
  4020 => (x"f2",x"c0",x"87",x"e4"),
  4021 => (x"f0",x"fc",x"c3",x"1e"),
  4022 => (x"87",x"da",x"fb",x"49"),
  4023 => (x"48",x"cd",x"eb",x"c1"),
  4024 => (x"1e",x"c0",x"50",x"c1"),
  4025 => (x"bf",x"cc",x"c4",x"c4"),
  4026 => (x"87",x"ca",x"fb",x"49"),
  4027 => (x"98",x"70",x"86",x"cc"),
  4028 => (x"c3",x"87",x"c4",x"05"),
  4029 => (x"c4",x"4b",x"fc",x"fc"),
  4030 => (x"48",x"bf",x"ea",x"d9"),
  4031 => (x"d9",x"c4",x"98",x"fd"),
  4032 => (x"e7",x"f6",x"58",x"ee"),
  4033 => (x"87",x"ee",x"e8",x"87"),
  4034 => (x"87",x"ce",x"f1",x"fd"),
  4035 => (x"ff",x"fd",x"49",x"c1"),
  4036 => (x"c8",x"c3",x"87",x"f5"),
  4037 => (x"c3",x"1e",x"c1",x"1e"),
  4038 => (x"f8",x"e8",x"49",x"ff"),
  4039 => (x"f8",x"48",x"73",x"87"),
  4040 => (x"87",x"ca",x"e8",x"8e"),
  4041 => (x"53",x"4f",x"4d",x"43"),
  4042 => (x"20",x"20",x"20",x"20"),
  4043 => (x"00",x"4d",x"41",x"52"),
  4044 => (x"48",x"43",x"52",x"41"),
  4045 => (x"20",x"31",x"45",x"49"),
  4046 => (x"00",x"46",x"44",x"48"),
  4047 => (x"20",x"4d",x"4f",x"52"),
  4048 => (x"64",x"61",x"6f",x"6c"),
  4049 => (x"20",x"67",x"6e",x"69"),
  4050 => (x"6c",x"69",x"61",x"66"),
  4051 => (x"00",x"2e",x"64",x"65"),
  4052 => (x"1e",x"1e",x"73",x"1e"),
  4053 => (x"fe",x"fd",x"49",x"c0"),
  4054 => (x"e7",x"e9",x"87",x"ed"),
  4055 => (x"fe",x"4b",x"70",x"87"),
  4056 => (x"73",x"87",x"ee",x"df"),
  4057 => (x"87",x"c8",x"05",x"9b"),
  4058 => (x"87",x"da",x"eb",x"fe"),
  4059 => (x"87",x"e5",x"d3",x"ff"),
  4060 => (x"ff",x"c1",x"49",x"6e"),
  4061 => (x"48",x"6e",x"99",x"ff"),
  4062 => (x"7e",x"70",x"80",x"c1"),
  4063 => (x"ff",x"05",x"99",x"71"),
  4064 => (x"e9",x"fd",x"87",x"d2"),
  4065 => (x"49",x"70",x"87",x"cf"),
  4066 => (x"87",x"d3",x"c6",x"fe"),
  4067 => (x"26",x"87",x"c5",x"ff"),
  4068 => (x"76",x"87",x"db",x"e6"),
  4069 => (x"0c",x"04",x"06",x"05"),
  4070 => (x"0a",x"83",x"0b",x"03"),
  4071 => (x"07",x"78",x"09",x"01"),
  4072 => (x"0e",x"f7",x"7e",x"fc"),
  4073 => (x"25",x"26",x"1e",x"16"),
  4074 => (x"3e",x"3d",x"36",x"2e"),
  4075 => (x"55",x"7b",x"45",x"46"),
  4076 => (x"ec",x"f0",x"66",x"ff"),
  4077 => (x"7c",x"ca",x"77",x"fd"),
  4078 => (x"1d",x"15",x"0d",x"ff"),
  4079 => (x"35",x"2c",x"2d",x"24"),
  4080 => (x"4d",x"44",x"43",x"3c"),
  4081 => (x"f1",x"5d",x"5b",x"54"),
  4082 => (x"75",x"6c",x"fa",x"e9"),
  4083 => (x"1c",x"14",x"84",x"7d"),
  4084 => (x"34",x"2b",x"23",x"1b"),
  4085 => (x"4b",x"42",x"3b",x"33"),
  4086 => (x"6b",x"5a",x"52",x"4c"),
  4087 => (x"12",x"79",x"74",x"73"),
  4088 => (x"21",x"22",x"1a",x"ff"),
  4089 => (x"3a",x"31",x"32",x"2a"),
  4090 => (x"59",x"4a",x"49",x"41"),
  4091 => (x"7a",x"72",x"69",x"f5"),
  4092 => (x"91",x"29",x"11",x"58"),
  4093 => (x"f4",x"f2",x"eb",x"94"),
  4094 => (x"00",x"da",x"71",x"70"),
  4095 => (x"f5",x"f2",x"eb",x"f4"),
  4096 => (x"0c",x"04",x"06",x"05"),
  4097 => (x"0a",x"83",x"0b",x"03"),
  4098 => (x"00",x"07",x"00",x"66"),
  4099 => (x"00",x"da",x"00",x"5a"),
  4100 => (x"08",x"94",x"80",x"00"),
  4101 => (x"00",x"07",x"80",x"05"),
  4102 => (x"00",x"01",x"80",x"02"),
  4103 => (x"00",x"09",x"80",x"03"),
  4104 => (x"00",x"78",x"80",x"04"),
  4105 => (x"08",x"91",x"80",x"01"),
  4106 => (x"00",x"00",x"00",x"26"),
  4107 => (x"00",x"00",x"00",x"1d"),
  4108 => (x"00",x"00",x"00",x"1c"),
  4109 => (x"00",x"00",x"00",x"25"),
  4110 => (x"00",x"00",x"00",x"1a"),
  4111 => (x"00",x"00",x"00",x"1b"),
  4112 => (x"00",x"00",x"00",x"24"),
  4113 => (x"00",x"00",x"01",x"12"),
  4114 => (x"00",x"00",x"00",x"2e"),
  4115 => (x"00",x"00",x"00",x"2d"),
  4116 => (x"00",x"00",x"00",x"23"),
  4117 => (x"00",x"00",x"00",x"36"),
  4118 => (x"00",x"00",x"00",x"21"),
  4119 => (x"00",x"00",x"00",x"2b"),
  4120 => (x"00",x"00",x"00",x"2c"),
  4121 => (x"00",x"00",x"00",x"22"),
  4122 => (x"00",x"6c",x"00",x"3d"),
  4123 => (x"00",x"00",x"00",x"35"),
  4124 => (x"00",x"00",x"00",x"34"),
  4125 => (x"00",x"75",x"00",x"3e"),
  4126 => (x"00",x"00",x"00",x"32"),
  4127 => (x"00",x"00",x"00",x"33"),
  4128 => (x"00",x"6b",x"00",x"3c"),
  4129 => (x"00",x"00",x"00",x"2a"),
  4130 => (x"00",x"7d",x"00",x"46"),
  4131 => (x"00",x"73",x"00",x"43"),
  4132 => (x"00",x"69",x"00",x"3b"),
  4133 => (x"00",x"ca",x"00",x"45"),
  4134 => (x"00",x"70",x"00",x"3a"),
  4135 => (x"00",x"72",x"00",x"42"),
  4136 => (x"00",x"74",x"00",x"44"),
  4137 => (x"00",x"00",x"00",x"31"),
  4138 => (x"00",x"78",x"00",x"55"),
  4139 => (x"00",x"7c",x"00",x"4d"),
  4140 => (x"00",x"7a",x"00",x"4b"),
  4141 => (x"00",x"7e",x"00",x"7b"),
  4142 => (x"00",x"71",x"00",x"49"),
  4143 => (x"00",x"84",x"00",x"4c"),
  4144 => (x"00",x"77",x"00",x"54"),
  4145 => (x"00",x"00",x"00",x"41"),
  4146 => (x"00",x"fc",x"00",x"61"),
  4147 => (x"00",x"7c",x"00",x"5b"),
  4148 => (x"00",x"00",x"00",x"52"),
  4149 => (x"00",x"78",x"00",x"f1"),
  4150 => (x"00",x"00",x"02",x"59"),
  4151 => (x"00",x"5d",x"00",x"0e"),
  4152 => (x"00",x"00",x"00",x"5d"),
  4153 => (x"00",x"79",x"00",x"4a"),
  4154 => (x"00",x"00",x"00",x"16"),
  4155 => (x"00",x"fc",x"00",x"76"),
  4156 => (x"00",x"0d",x"04",x"14"),
  4157 => (x"00",x"00",x"00",x"1e"),
  4158 => (x"00",x"00",x"00",x"29"),
  4159 => (x"00",x"00",x"00",x"11"),
  4160 => (x"00",x"00",x"00",x"15"),
  4161 => (x"00",x"00",x"40",x"00"),
  4162 => (x"00",x"00",x"41",x"10"),
  4163 => (x"00",x"00",x"41",x"a5"),
  4164 => (x"3b",x"63",x"72",x"41"),
  4165 => (x"3b",x"4d",x"4f",x"52"),
  4166 => (x"2c",x"55",x"30",x"53"),
  4167 => (x"2c",x"46",x"44",x"41"),
  4168 => (x"70",x"6f",x"6c",x"46"),
  4169 => (x"31",x"20",x"79",x"70"),
  4170 => (x"31",x"53",x"3b",x"3a"),
  4171 => (x"44",x"41",x"2c",x"55"),
  4172 => (x"6c",x"46",x"2c",x"46"),
  4173 => (x"79",x"70",x"70",x"6f"),
  4174 => (x"3b",x"3a",x"32",x"20"),
  4175 => (x"2c",x"55",x"32",x"53"),
  4176 => (x"2c",x"46",x"44",x"48"),
  4177 => (x"64",x"72",x"61",x"48"),
  4178 => (x"73",x"69",x"64",x"20"),
  4179 => (x"3a",x"31",x"20",x"6b"),
  4180 => (x"55",x"33",x"53",x"3b"),
  4181 => (x"46",x"44",x"48",x"2c"),
  4182 => (x"72",x"61",x"48",x"2c"),
  4183 => (x"69",x"64",x"20",x"64"),
  4184 => (x"32",x"20",x"6b",x"73"),
  4185 => (x"52",x"53",x"3b",x"3a"),
  4186 => (x"41",x"52",x"2c",x"55"),
  4187 => (x"6f",x"4c",x"2c",x"4d"),
  4188 => (x"43",x"20",x"64",x"61"),
  4189 => (x"20",x"53",x"4f",x"4d"),
  4190 => (x"3a",x"4d",x"41",x"52"),
  4191 => (x"55",x"53",x"53",x"3b"),
  4192 => (x"4d",x"41",x"52",x"2c"),
  4193 => (x"76",x"61",x"53",x"2c"),
  4194 => (x"4d",x"43",x"20",x"65"),
  4195 => (x"52",x"20",x"53",x"4f"),
  4196 => (x"3b",x"3a",x"4d",x"41"),
  4197 => (x"52",x"2c",x"31",x"54"),
  4198 => (x"74",x"65",x"73",x"65"),
  4199 => (x"76",x"2c",x"56",x"3b"),
  4200 => (x"2e",x"30",x"2e",x"31"),
  4201 => (x"53",x"49",x"52",x"00"),
  4202 => (x"20",x"53",x"4f",x"43"),
  4203 => (x"4d",x"4f",x"52",x"20"),
  4204 => (x"4d",x"4f",x"52",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

